// This is the unpowered netlist.
module tt_um_hsc_tdc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net16;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire tdc_inst_capt_out_0 ;
 wire tdc_inst_capt_out_10 ;
 wire tdc_inst_capt_out_11 ;
 wire tdc_inst_capt_out_12 ;
 wire tdc_inst_capt_out_13 ;
 wire tdc_inst_capt_out_14 ;
 wire tdc_inst_capt_out_15 ;
 wire tdc_inst_capt_out_16 ;
 wire tdc_inst_capt_out_17 ;
 wire tdc_inst_capt_out_18 ;
 wire tdc_inst_capt_out_19 ;
 wire tdc_inst_capt_out_1 ;
 wire tdc_inst_capt_out_20 ;
 wire tdc_inst_capt_out_21 ;
 wire tdc_inst_capt_out_22 ;
 wire tdc_inst_capt_out_23 ;
 wire tdc_inst_capt_out_24 ;
 wire tdc_inst_capt_out_25 ;
 wire tdc_inst_capt_out_26 ;
 wire tdc_inst_capt_out_27 ;
 wire tdc_inst_capt_out_28 ;
 wire tdc_inst_capt_out_29 ;
 wire tdc_inst_capt_out_2 ;
 wire tdc_inst_capt_out_30 ;
 wire tdc_inst_capt_out_31 ;
 wire tdc_inst_capt_out_32 ;
 wire tdc_inst_capt_out_33 ;
 wire tdc_inst_capt_out_34 ;
 wire tdc_inst_capt_out_35 ;
 wire tdc_inst_capt_out_36 ;
 wire tdc_inst_capt_out_37 ;
 wire tdc_inst_capt_out_38 ;
 wire tdc_inst_capt_out_39 ;
 wire tdc_inst_capt_out_3 ;
 wire tdc_inst_capt_out_40 ;
 wire tdc_inst_capt_out_41 ;
 wire tdc_inst_capt_out_42 ;
 wire tdc_inst_capt_out_43 ;
 wire tdc_inst_capt_out_44 ;
 wire tdc_inst_capt_out_45 ;
 wire tdc_inst_capt_out_46 ;
 wire tdc_inst_capt_out_47 ;
 wire tdc_inst_capt_out_48 ;
 wire tdc_inst_capt_out_49 ;
 wire tdc_inst_capt_out_4 ;
 wire tdc_inst_capt_out_50 ;
 wire tdc_inst_capt_out_51 ;
 wire tdc_inst_capt_out_52 ;
 wire tdc_inst_capt_out_53 ;
 wire tdc_inst_capt_out_54 ;
 wire tdc_inst_capt_out_55 ;
 wire tdc_inst_capt_out_56 ;
 wire tdc_inst_capt_out_57 ;
 wire tdc_inst_capt_out_58 ;
 wire tdc_inst_capt_out_59 ;
 wire tdc_inst_capt_out_5 ;
 wire tdc_inst_capt_out_60 ;
 wire tdc_inst_capt_out_61 ;
 wire tdc_inst_capt_out_62 ;
 wire tdc_inst_capt_out_63 ;
 wire tdc_inst_capt_out_6 ;
 wire tdc_inst_capt_out_7 ;
 wire tdc_inst_capt_out_8 ;
 wire tdc_inst_capt_out_9 ;
 wire tdc_inst_capt_reg_r_1_0 ;
 wire tdc_inst_capt_reg_r_1_10 ;
 wire tdc_inst_capt_reg_r_1_11 ;
 wire tdc_inst_capt_reg_r_1_12 ;
 wire tdc_inst_capt_reg_r_1_13 ;
 wire tdc_inst_capt_reg_r_1_14 ;
 wire tdc_inst_capt_reg_r_1_15 ;
 wire tdc_inst_capt_reg_r_1_16 ;
 wire tdc_inst_capt_reg_r_1_17 ;
 wire tdc_inst_capt_reg_r_1_18 ;
 wire tdc_inst_capt_reg_r_1_19 ;
 wire tdc_inst_capt_reg_r_1_1 ;
 wire tdc_inst_capt_reg_r_1_20 ;
 wire tdc_inst_capt_reg_r_1_21 ;
 wire tdc_inst_capt_reg_r_1_22 ;
 wire tdc_inst_capt_reg_r_1_23 ;
 wire tdc_inst_capt_reg_r_1_24 ;
 wire tdc_inst_capt_reg_r_1_25 ;
 wire tdc_inst_capt_reg_r_1_26 ;
 wire tdc_inst_capt_reg_r_1_27 ;
 wire tdc_inst_capt_reg_r_1_28 ;
 wire tdc_inst_capt_reg_r_1_29 ;
 wire tdc_inst_capt_reg_r_1_2 ;
 wire tdc_inst_capt_reg_r_1_30 ;
 wire tdc_inst_capt_reg_r_1_31 ;
 wire tdc_inst_capt_reg_r_1_32 ;
 wire tdc_inst_capt_reg_r_1_33 ;
 wire tdc_inst_capt_reg_r_1_34 ;
 wire tdc_inst_capt_reg_r_1_35 ;
 wire tdc_inst_capt_reg_r_1_36 ;
 wire tdc_inst_capt_reg_r_1_37 ;
 wire tdc_inst_capt_reg_r_1_38 ;
 wire tdc_inst_capt_reg_r_1_39 ;
 wire tdc_inst_capt_reg_r_1_3 ;
 wire tdc_inst_capt_reg_r_1_40 ;
 wire tdc_inst_capt_reg_r_1_41 ;
 wire tdc_inst_capt_reg_r_1_42 ;
 wire tdc_inst_capt_reg_r_1_43 ;
 wire tdc_inst_capt_reg_r_1_44 ;
 wire tdc_inst_capt_reg_r_1_45 ;
 wire tdc_inst_capt_reg_r_1_46 ;
 wire tdc_inst_capt_reg_r_1_47 ;
 wire tdc_inst_capt_reg_r_1_48 ;
 wire tdc_inst_capt_reg_r_1_49 ;
 wire tdc_inst_capt_reg_r_1_4 ;
 wire tdc_inst_capt_reg_r_1_50 ;
 wire tdc_inst_capt_reg_r_1_51 ;
 wire tdc_inst_capt_reg_r_1_52 ;
 wire tdc_inst_capt_reg_r_1_53 ;
 wire tdc_inst_capt_reg_r_1_54 ;
 wire tdc_inst_capt_reg_r_1_55 ;
 wire tdc_inst_capt_reg_r_1_56 ;
 wire tdc_inst_capt_reg_r_1_57 ;
 wire tdc_inst_capt_reg_r_1_58 ;
 wire tdc_inst_capt_reg_r_1_59 ;
 wire tdc_inst_capt_reg_r_1_5 ;
 wire tdc_inst_capt_reg_r_1_60 ;
 wire tdc_inst_capt_reg_r_1_61 ;
 wire tdc_inst_capt_reg_r_1_62 ;
 wire tdc_inst_capt_reg_r_1_63 ;
 wire tdc_inst_capt_reg_r_1_6 ;
 wire tdc_inst_capt_reg_r_1_7 ;
 wire tdc_inst_capt_reg_r_1_8 ;
 wire tdc_inst_capt_reg_r_1_9 ;
 wire tdc_inst_dl_capt_D_0 ;
 wire tdc_inst_dl_capt_D_10 ;
 wire tdc_inst_dl_capt_D_11 ;
 wire tdc_inst_dl_capt_D_12 ;
 wire tdc_inst_dl_capt_D_13 ;
 wire tdc_inst_dl_capt_D_14 ;
 wire tdc_inst_dl_capt_D_15 ;
 wire tdc_inst_dl_capt_D_16 ;
 wire tdc_inst_dl_capt_D_17 ;
 wire tdc_inst_dl_capt_D_18 ;
 wire tdc_inst_dl_capt_D_19 ;
 wire tdc_inst_dl_capt_D_1 ;
 wire tdc_inst_dl_capt_D_20 ;
 wire tdc_inst_dl_capt_D_21 ;
 wire tdc_inst_dl_capt_D_22 ;
 wire tdc_inst_dl_capt_D_23 ;
 wire tdc_inst_dl_capt_D_24 ;
 wire tdc_inst_dl_capt_D_25 ;
 wire tdc_inst_dl_capt_D_26 ;
 wire tdc_inst_dl_capt_D_27 ;
 wire tdc_inst_dl_capt_D_28 ;
 wire tdc_inst_dl_capt_D_29 ;
 wire tdc_inst_dl_capt_D_2 ;
 wire tdc_inst_dl_capt_D_30 ;
 wire tdc_inst_dl_capt_D_31 ;
 wire tdc_inst_dl_capt_D_32 ;
 wire tdc_inst_dl_capt_D_33 ;
 wire tdc_inst_dl_capt_D_34 ;
 wire tdc_inst_dl_capt_D_35 ;
 wire tdc_inst_dl_capt_D_36 ;
 wire tdc_inst_dl_capt_D_37 ;
 wire tdc_inst_dl_capt_D_38 ;
 wire tdc_inst_dl_capt_D_39 ;
 wire tdc_inst_dl_capt_D_3 ;
 wire tdc_inst_dl_capt_D_40 ;
 wire tdc_inst_dl_capt_D_41 ;
 wire tdc_inst_dl_capt_D_42 ;
 wire tdc_inst_dl_capt_D_43 ;
 wire tdc_inst_dl_capt_D_44 ;
 wire tdc_inst_dl_capt_D_45 ;
 wire tdc_inst_dl_capt_D_46 ;
 wire tdc_inst_dl_capt_D_47 ;
 wire tdc_inst_dl_capt_D_48 ;
 wire tdc_inst_dl_capt_D_49 ;
 wire tdc_inst_dl_capt_D_4 ;
 wire tdc_inst_dl_capt_D_50 ;
 wire tdc_inst_dl_capt_D_51 ;
 wire tdc_inst_dl_capt_D_52 ;
 wire tdc_inst_dl_capt_D_53 ;
 wire tdc_inst_dl_capt_D_54 ;
 wire tdc_inst_dl_capt_D_55 ;
 wire tdc_inst_dl_capt_D_56 ;
 wire tdc_inst_dl_capt_D_57 ;
 wire tdc_inst_dl_capt_D_58 ;
 wire tdc_inst_dl_capt_D_59 ;
 wire tdc_inst_dl_capt_D_5 ;
 wire tdc_inst_dl_capt_D_60 ;
 wire tdc_inst_dl_capt_D_61 ;
 wire tdc_inst_dl_capt_D_62 ;
 wire tdc_inst_dl_capt_D_63 ;
 wire tdc_inst_dl_capt_D_6 ;
 wire tdc_inst_dl_capt_D_7 ;
 wire tdc_inst_dl_capt_D_8 ;
 wire tdc_inst_dl_capt_D_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_0 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_10 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_11 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_12 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_13 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_14 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_15 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_16 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_17 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_18 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_19 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_1 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_20 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_21 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_22 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_23 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_24 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_25 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_26 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_27 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_28 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_29 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_2 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_30 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_31 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_32 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_33 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_34 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_35 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_36 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_37 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_38 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_39 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_3 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_40 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_41 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_42 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_43 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_44 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_45 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_46 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_47 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_48 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_49 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_4 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_50 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_51 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_52 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_53 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_54 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_55 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_56 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_57 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_58 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_59 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_5 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_60 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_61 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_62 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_63 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_6 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_7 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_8 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_9 ;
 wire tdc_inst_dl_inst_dl_genblk_keep_co ;
 wire tdc_inst_pg_pg_r_out ;
 wire [1:0] clknet_0_ui_in;
 wire [1:0] clknet_4_0_0_ui_in;
 wire [1:0] clknet_4_10_0_ui_in;
 wire [1:0] clknet_4_11_0_ui_in;
 wire [1:0] clknet_4_12_0_ui_in;
 wire [1:0] clknet_4_13_0_ui_in;
 wire [1:0] clknet_4_14_0_ui_in;
 wire [1:0] clknet_4_15_0_ui_in;
 wire [1:0] clknet_4_1_0_ui_in;
 wire [1:0] clknet_4_2_0_ui_in;
 wire [1:0] clknet_4_3_0_ui_in;
 wire [1:0] clknet_4_4_0_ui_in;
 wire [1:0] clknet_4_5_0_ui_in;
 wire [1:0] clknet_4_6_0_ui_in;
 wire [1:0] clknet_4_7_0_ui_in;
 wire [1:0] clknet_4_8_0_ui_in;
 wire [1:0] clknet_4_9_0_ui_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__mux2_4 _0643_ (.A0(net6),
    .A1(tdc_inst_pg_pg_r_out ),
    .S(net4),
    .X(_0072_));
 sky130_fd_sc_hd__buf_6 _0644_ (.A(_0072_),
    .X(tdc_inst_dl_inst_dl_genblk_dl_c_0 ));
 sky130_fd_sc_hd__buf_2 _0645_ (.A(net2),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(net5),
    .A1(net6),
    .S(net3),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_4 _0647_ (.A(net16),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0648_ (.A0(tdc_inst_pg_pg_r_out ),
    .A1(_0074_),
    .S(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _0649_ (.A(_0073_),
    .B(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(_0077_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _0651_ (.A0(tdc_inst_capt_reg_r_1_0 ),
    .A1(tdc_inst_capt_out_0 ),
    .S(_0075_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _0652_ (.A(_0073_),
    .B(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _0653_ (.A(_0079_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0654_ (.A0(tdc_inst_capt_reg_r_1_1 ),
    .A1(tdc_inst_capt_out_1 ),
    .S(_0075_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _0655_ (.A(_0073_),
    .B(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _0656_ (.A(_0081_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_2 _0657_ (.A(net2),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(tdc_inst_capt_reg_r_1_2 ),
    .A1(tdc_inst_capt_out_2 ),
    .S(_0075_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _0659_ (.A(_0082_),
    .B(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0084_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0661_ (.A0(tdc_inst_capt_reg_r_1_3 ),
    .A1(tdc_inst_capt_out_3 ),
    .S(_0075_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _0662_ (.A(_0082_),
    .B(_0085_),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _0663_ (.A(_0086_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(tdc_inst_capt_reg_r_1_4 ),
    .A1(tdc_inst_capt_out_4 ),
    .S(_0075_),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _0665_ (.A(_0082_),
    .B(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(_0088_),
    .X(_0005_));
 sky130_fd_sc_hd__buf_4 _0667_ (.A(net11),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_4 _0668_ (.A(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0669_ (.A0(tdc_inst_capt_reg_r_1_5 ),
    .A1(tdc_inst_capt_out_5 ),
    .S(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _0670_ (.A(_0082_),
    .B(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _0671_ (.A(_0092_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(tdc_inst_capt_reg_r_1_6 ),
    .A1(tdc_inst_capt_out_6 ),
    .S(_0090_),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _0673_ (.A(_0082_),
    .B(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _0674_ (.A(_0094_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0675_ (.A0(tdc_inst_capt_reg_r_1_7 ),
    .A1(tdc_inst_capt_out_7 ),
    .S(_0090_),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _0676_ (.A(_0082_),
    .B(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _0677_ (.A(_0096_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(tdc_inst_capt_reg_r_1_8 ),
    .A1(tdc_inst_capt_out_8 ),
    .S(_0090_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _0679_ (.A(_0082_),
    .B(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(_0098_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0681_ (.A0(tdc_inst_capt_reg_r_1_9 ),
    .A1(tdc_inst_capt_out_9 ),
    .S(_0090_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _0682_ (.A(_0082_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0683_ (.A(_0100_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(tdc_inst_capt_reg_r_1_10 ),
    .A1(tdc_inst_capt_out_10 ),
    .S(_0090_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _0685_ (.A(_0082_),
    .B(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _0686_ (.A(_0102_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(tdc_inst_capt_reg_r_1_11 ),
    .A1(tdc_inst_capt_out_11 ),
    .S(_0090_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _0688_ (.A(_0082_),
    .B(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0689_ (.A(_0104_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_2 _0690_ (.A(net2),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(tdc_inst_capt_reg_r_1_12 ),
    .A1(tdc_inst_capt_out_12 ),
    .S(_0090_),
    .X(_0106_));
 sky130_fd_sc_hd__and2_1 _0692_ (.A(_0105_),
    .B(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0693_ (.A(_0107_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(tdc_inst_capt_reg_r_1_13 ),
    .A1(tdc_inst_capt_out_13 ),
    .S(_0090_),
    .X(_0108_));
 sky130_fd_sc_hd__and2_1 _0695_ (.A(_0105_),
    .B(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0696_ (.A(_0109_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(tdc_inst_capt_reg_r_1_14 ),
    .A1(tdc_inst_capt_out_14 ),
    .S(_0090_),
    .X(_0110_));
 sky130_fd_sc_hd__and2_1 _0698_ (.A(_0105_),
    .B(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _0699_ (.A(_0111_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_4 _0700_ (.A(net14),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0701_ (.A0(tdc_inst_capt_reg_r_1_15 ),
    .A1(tdc_inst_capt_out_15 ),
    .S(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__and2_1 _0702_ (.A(_0105_),
    .B(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0114_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(tdc_inst_capt_reg_r_1_16 ),
    .A1(tdc_inst_capt_out_16 ),
    .S(_0112_),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _0705_ (.A(_0105_),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0706_ (.A(_0116_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(tdc_inst_capt_reg_r_1_17 ),
    .A1(tdc_inst_capt_out_17 ),
    .S(_0112_),
    .X(_0117_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(_0105_),
    .B(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0118_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(tdc_inst_capt_reg_r_1_18 ),
    .A1(tdc_inst_capt_out_18 ),
    .S(_0112_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(_0105_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0120_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(tdc_inst_capt_reg_r_1_19 ),
    .A1(tdc_inst_capt_out_19 ),
    .S(_0112_),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _0714_ (.A(_0105_),
    .B(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _0715_ (.A(_0122_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(tdc_inst_capt_reg_r_1_20 ),
    .A1(tdc_inst_capt_out_20 ),
    .S(_0112_),
    .X(_0123_));
 sky130_fd_sc_hd__and2_1 _0717_ (.A(_0105_),
    .B(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0718_ (.A(_0124_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(tdc_inst_capt_reg_r_1_21 ),
    .A1(tdc_inst_capt_out_21 ),
    .S(_0112_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _0720_ (.A(_0105_),
    .B(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0721_ (.A(_0126_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_2 _0722_ (.A(net2),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(tdc_inst_capt_reg_r_1_22 ),
    .A1(tdc_inst_capt_out_22 ),
    .S(_0112_),
    .X(_0128_));
 sky130_fd_sc_hd__and2_1 _0724_ (.A(_0127_),
    .B(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _0725_ (.A(_0129_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(tdc_inst_capt_reg_r_1_23 ),
    .A1(tdc_inst_capt_out_23 ),
    .S(_0112_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(_0127_),
    .B(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _0728_ (.A(_0131_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(tdc_inst_capt_reg_r_1_24 ),
    .A1(tdc_inst_capt_out_24 ),
    .S(_0112_),
    .X(_0132_));
 sky130_fd_sc_hd__and2_1 _0730_ (.A(_0127_),
    .B(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _0731_ (.A(_0133_),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_4 _0732_ (.A(net9),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0733_ (.A0(tdc_inst_capt_reg_r_1_25 ),
    .A1(tdc_inst_capt_out_25 ),
    .S(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _0734_ (.A(_0127_),
    .B(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0136_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(tdc_inst_capt_reg_r_1_26 ),
    .A1(tdc_inst_capt_out_26 ),
    .S(_0134_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_1 _0737_ (.A(_0127_),
    .B(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0738_ (.A(_0138_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0739_ (.A0(tdc_inst_capt_reg_r_1_27 ),
    .A1(tdc_inst_capt_out_27 ),
    .S(_0134_),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _0740_ (.A(_0127_),
    .B(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _0741_ (.A(_0140_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(tdc_inst_capt_reg_r_1_28 ),
    .A1(tdc_inst_capt_out_28 ),
    .S(_0134_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _0743_ (.A(_0127_),
    .B(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0744_ (.A(_0142_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0745_ (.A0(tdc_inst_capt_reg_r_1_29 ),
    .A1(tdc_inst_capt_out_29 ),
    .S(_0134_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _0746_ (.A(_0127_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0144_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(tdc_inst_capt_reg_r_1_30 ),
    .A1(tdc_inst_capt_out_30 ),
    .S(_0134_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _0749_ (.A(_0127_),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0750_ (.A(_0146_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0751_ (.A0(tdc_inst_capt_reg_r_1_31 ),
    .A1(tdc_inst_capt_out_31 ),
    .S(_0134_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_1 _0752_ (.A(_0127_),
    .B(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0148_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_2 _0754_ (.A(net2),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(tdc_inst_capt_reg_r_1_32 ),
    .A1(tdc_inst_capt_out_32 ),
    .S(_0134_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_1 _0756_ (.A(_0149_),
    .B(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0151_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(tdc_inst_capt_reg_r_1_33 ),
    .A1(tdc_inst_capt_out_33 ),
    .S(_0134_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_1 _0759_ (.A(_0149_),
    .B(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _0760_ (.A(_0153_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(tdc_inst_capt_reg_r_1_34 ),
    .A1(tdc_inst_capt_out_34 ),
    .S(_0134_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_1 _0762_ (.A(_0149_),
    .B(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0763_ (.A(_0155_),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_4 _0764_ (.A(net11),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(tdc_inst_capt_reg_r_1_35 ),
    .A1(tdc_inst_capt_out_35 ),
    .S(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _0766_ (.A(_0149_),
    .B(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0767_ (.A(_0158_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(tdc_inst_capt_reg_r_1_36 ),
    .A1(tdc_inst_capt_out_36 ),
    .S(_0156_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _0769_ (.A(_0149_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(_0160_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(tdc_inst_capt_reg_r_1_37 ),
    .A1(tdc_inst_capt_out_37 ),
    .S(_0156_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _0772_ (.A(_0149_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _0773_ (.A(_0162_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0774_ (.A0(tdc_inst_capt_reg_r_1_38 ),
    .A1(tdc_inst_capt_out_38 ),
    .S(_0156_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(_0149_),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0776_ (.A(_0164_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(tdc_inst_capt_reg_r_1_39 ),
    .A1(tdc_inst_capt_out_39 ),
    .S(_0156_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_1 _0778_ (.A(_0149_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0779_ (.A(_0166_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(tdc_inst_capt_reg_r_1_40 ),
    .A1(tdc_inst_capt_out_40 ),
    .S(_0156_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _0781_ (.A(_0149_),
    .B(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0782_ (.A(_0168_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(tdc_inst_capt_reg_r_1_41 ),
    .A1(tdc_inst_capt_out_41 ),
    .S(_0156_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _0784_ (.A(_0149_),
    .B(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0785_ (.A(_0170_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_2 _0786_ (.A(net2),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(tdc_inst_capt_reg_r_1_42 ),
    .A1(tdc_inst_capt_out_42 ),
    .S(_0156_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _0788_ (.A(_0171_),
    .B(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _0789_ (.A(_0173_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(tdc_inst_capt_reg_r_1_43 ),
    .A1(tdc_inst_capt_out_43 ),
    .S(_0156_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _0791_ (.A(_0171_),
    .B(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _0792_ (.A(_0175_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(tdc_inst_capt_reg_r_1_44 ),
    .A1(tdc_inst_capt_out_44 ),
    .S(_0156_),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _0794_ (.A(_0171_),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_1 _0795_ (.A(_0177_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _0796_ (.A(net11),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(tdc_inst_capt_reg_r_1_45 ),
    .A1(tdc_inst_capt_out_45 ),
    .S(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_1 _0798_ (.A(_0171_),
    .B(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _0799_ (.A(_0180_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(tdc_inst_capt_reg_r_1_46 ),
    .A1(tdc_inst_capt_out_46 ),
    .S(_0178_),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _0801_ (.A(_0171_),
    .B(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(_0182_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0803_ (.A0(tdc_inst_capt_reg_r_1_47 ),
    .A1(tdc_inst_capt_out_47 ),
    .S(_0178_),
    .X(_0183_));
 sky130_fd_sc_hd__and2_1 _0804_ (.A(_0171_),
    .B(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0805_ (.A(_0184_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(tdc_inst_capt_reg_r_1_48 ),
    .A1(tdc_inst_capt_out_48 ),
    .S(_0178_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _0807_ (.A(_0171_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0808_ (.A(_0186_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(tdc_inst_capt_reg_r_1_49 ),
    .A1(tdc_inst_capt_out_49 ),
    .S(_0178_),
    .X(_0187_));
 sky130_fd_sc_hd__and2_1 _0810_ (.A(_0171_),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0188_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0812_ (.A0(tdc_inst_capt_reg_r_1_50 ),
    .A1(tdc_inst_capt_out_50 ),
    .S(_0178_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _0813_ (.A(_0171_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _0814_ (.A(_0190_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0815_ (.A0(tdc_inst_capt_reg_r_1_51 ),
    .A1(tdc_inst_capt_out_51 ),
    .S(_0178_),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _0816_ (.A(_0171_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0817_ (.A(_0192_),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_2 _0818_ (.A(net2),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _0819_ (.A0(tdc_inst_capt_reg_r_1_52 ),
    .A1(tdc_inst_capt_out_52 ),
    .S(_0178_),
    .X(_0194_));
 sky130_fd_sc_hd__and2_1 _0820_ (.A(_0193_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _0821_ (.A(_0195_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0822_ (.A0(tdc_inst_capt_reg_r_1_53 ),
    .A1(tdc_inst_capt_out_53 ),
    .S(_0178_),
    .X(_0196_));
 sky130_fd_sc_hd__and2_1 _0823_ (.A(_0193_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0197_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(tdc_inst_capt_reg_r_1_54 ),
    .A1(tdc_inst_capt_out_54 ),
    .S(_0178_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_1 _0826_ (.A(_0193_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _0827_ (.A(_0199_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(tdc_inst_capt_reg_r_1_55 ),
    .A1(tdc_inst_capt_out_55 ),
    .S(_0089_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _0829_ (.A(_0193_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _0830_ (.A(_0201_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(tdc_inst_capt_reg_r_1_56 ),
    .A1(tdc_inst_capt_out_56 ),
    .S(_0089_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _0832_ (.A(_0193_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _0833_ (.A(_0203_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0834_ (.A0(tdc_inst_capt_reg_r_1_57 ),
    .A1(tdc_inst_capt_out_57 ),
    .S(_0089_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _0835_ (.A(_0193_),
    .B(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(_0205_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(tdc_inst_capt_reg_r_1_58 ),
    .A1(tdc_inst_capt_out_58 ),
    .S(_0089_),
    .X(_0206_));
 sky130_fd_sc_hd__and2_1 _0838_ (.A(_0193_),
    .B(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _0839_ (.A(_0207_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(tdc_inst_capt_reg_r_1_59 ),
    .A1(tdc_inst_capt_out_59 ),
    .S(_0089_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_1 _0841_ (.A(_0193_),
    .B(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _0842_ (.A(_0209_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0843_ (.A0(tdc_inst_capt_reg_r_1_60 ),
    .A1(tdc_inst_capt_out_60 ),
    .S(_0089_),
    .X(_0210_));
 sky130_fd_sc_hd__and2_1 _0844_ (.A(_0193_),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _0845_ (.A(_0211_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(tdc_inst_capt_reg_r_1_61 ),
    .A1(tdc_inst_capt_out_61 ),
    .S(_0089_),
    .X(_0212_));
 sky130_fd_sc_hd__and2_1 _0847_ (.A(_0193_),
    .B(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0213_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(tdc_inst_capt_reg_r_1_62 ),
    .A1(tdc_inst_capt_out_62 ),
    .S(_0089_),
    .X(_0214_));
 sky130_fd_sc_hd__and2_1 _0850_ (.A(net2),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_1 _0851_ (.A(_0215_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(tdc_inst_capt_reg_r_1_63 ),
    .A1(tdc_inst_capt_out_63 ),
    .S(_0089_),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(net2),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _0854_ (.A(_0217_),
    .X(_0064_));
 sky130_fd_sc_hd__buf_2 _0855_ (.A(_0075_),
    .X(_0218_));
 sky130_fd_sc_hd__inv_2 _0856_ (.A(tdc_inst_capt_reg_r_1_59 ),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(tdc_inst_capt_reg_r_1_40 ),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _0858_ (.A(tdc_inst_capt_reg_r_1_57 ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0859_ (.A(tdc_inst_capt_reg_r_1_53 ),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _0860_ (.A(tdc_inst_capt_reg_r_1_49 ),
    .Y(_0223_));
 sky130_fd_sc_hd__or2_1 _0861_ (.A(tdc_inst_capt_reg_r_1_60 ),
    .B(tdc_inst_capt_reg_r_1_3 ),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _0862_ (.A(tdc_inst_capt_reg_r_1_60 ),
    .B(tdc_inst_capt_reg_r_1_3 ),
    .Y(_0225_));
 sky130_fd_sc_hd__nand2_1 _0863_ (.A(_0224_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__xor2_1 _0864_ (.A(tdc_inst_capt_reg_r_1_63 ),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(tdc_inst_capt_reg_r_1_9 ),
    .Y(_0228_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(tdc_inst_capt_reg_r_1_37 ),
    .B(tdc_inst_capt_reg_r_1_35 ),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(tdc_inst_capt_reg_r_1_37 ),
    .B(tdc_inst_capt_reg_r_1_35 ),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _0868_ (.A(_0229_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__xor2_1 _0869_ (.A(tdc_inst_capt_reg_r_1_41 ),
    .B(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__xnor2_1 _0870_ (.A(_0228_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__xor2_1 _0871_ (.A(_0227_),
    .B(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__xor2_1 _0872_ (.A(tdc_inst_capt_reg_r_1_27 ),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__xnor2_1 _0873_ (.A(tdc_inst_capt_reg_r_1_8 ),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _0874_ (.A(tdc_inst_capt_reg_r_1_36 ),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _0875_ (.A(tdc_inst_capt_reg_r_1_25 ),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(tdc_inst_capt_reg_r_1_21 ),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _0877_ (.A(tdc_inst_capt_reg_r_1_14 ),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _0878_ (.A(tdc_inst_capt_reg_r_1_18 ),
    .Y(_0241_));
 sky130_fd_sc_hd__xor2_1 _0879_ (.A(tdc_inst_capt_reg_r_1_16 ),
    .B(tdc_inst_capt_reg_r_1_7 ),
    .X(_0242_));
 sky130_fd_sc_hd__xnor2_1 _0880_ (.A(tdc_inst_capt_reg_r_1_22 ),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_1 _0881_ (.A(_0241_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__xnor2_1 _0882_ (.A(_0240_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__xnor2_1 _0883_ (.A(_0239_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__xnor2_1 _0884_ (.A(_0238_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__xnor2_1 _0885_ (.A(_0237_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__xor2_1 _0886_ (.A(_0236_),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(tdc_inst_capt_reg_r_1_46 ),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _0888_ (.A(tdc_inst_capt_reg_r_1_46 ),
    .B(_0249_),
    .Y(_0251_));
 sky130_fd_sc_hd__nand2_1 _0889_ (.A(_0250_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__xnor2_2 _0890_ (.A(_0223_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _0891_ (.A(tdc_inst_capt_reg_r_1_33 ),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _0892_ (.A(tdc_inst_capt_reg_r_1_31 ),
    .Y(_0255_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(tdc_inst_capt_reg_r_1_10 ),
    .B(tdc_inst_capt_reg_r_1_6 ),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_2 _0894_ (.A(tdc_inst_capt_reg_r_1_10 ),
    .B(tdc_inst_capt_reg_r_1_6 ),
    .Y(_0257_));
 sky130_fd_sc_hd__a21o_1 _0895_ (.A1(_0256_),
    .A2(_0257_),
    .B1(tdc_inst_capt_reg_r_1_12 ),
    .X(_0258_));
 sky130_fd_sc_hd__nand3_2 _0896_ (.A(tdc_inst_capt_reg_r_1_12 ),
    .B(_0256_),
    .C(_0257_),
    .Y(_0259_));
 sky130_fd_sc_hd__nand2_1 _0897_ (.A(_0258_),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _0898_ (.A(tdc_inst_capt_reg_r_1_20 ),
    .Y(_0261_));
 sky130_fd_sc_hd__xor2_1 _0899_ (.A(tdc_inst_capt_reg_r_1_15 ),
    .B(tdc_inst_capt_reg_r_1_0 ),
    .X(_0262_));
 sky130_fd_sc_hd__xnor2_1 _0900_ (.A(tdc_inst_capt_reg_r_1_11 ),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__xnor2_1 _0901_ (.A(_0261_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand2_1 _0902_ (.A(_0260_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__or2_1 _0903_ (.A(_0260_),
    .B(_0264_),
    .X(_0266_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(_0265_),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__inv_2 _0905_ (.A(tdc_inst_capt_reg_r_1_17 ),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _0906_ (.A(tdc_inst_capt_reg_r_1_24 ),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _0907_ (.A(tdc_inst_capt_reg_r_1_5 ),
    .Y(_0270_));
 sky130_fd_sc_hd__xor2_1 _0908_ (.A(tdc_inst_capt_reg_r_1_26 ),
    .B(tdc_inst_capt_reg_r_1_23 ),
    .X(_0271_));
 sky130_fd_sc_hd__xnor2_1 _0909_ (.A(tdc_inst_capt_reg_r_1_19 ),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__xnor2_1 _0910_ (.A(_0270_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__xnor2_1 _0911_ (.A(_0269_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__xnor2_1 _0912_ (.A(_0268_),
    .B(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__xor2_1 _0913_ (.A(_0267_),
    .B(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_1 _0914_ (.A(_0255_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_1 _0915_ (.A(_0255_),
    .B(_0276_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _0916_ (.A(_0277_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__xnor2_2 _0917_ (.A(_0254_),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(tdc_inst_capt_reg_r_1_13 ),
    .Y(_0281_));
 sky130_fd_sc_hd__or2_1 _0919_ (.A(tdc_inst_capt_reg_r_1_32 ),
    .B(tdc_inst_capt_reg_r_1_30 ),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _0920_ (.A(tdc_inst_capt_reg_r_1_32 ),
    .B(tdc_inst_capt_reg_r_1_30 ),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_2 _0921_ (.A(_0282_),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__xor2_4 _0922_ (.A(tdc_inst_capt_reg_r_1_28 ),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _0923_ (.A(tdc_inst_capt_reg_r_1_39 ),
    .Y(_0286_));
 sky130_fd_sc_hd__xor2_2 _0924_ (.A(tdc_inst_capt_reg_r_1_42 ),
    .B(tdc_inst_capt_reg_r_1_38 ),
    .X(_0287_));
 sky130_fd_sc_hd__xnor2_2 _0925_ (.A(tdc_inst_capt_reg_r_1_34 ),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__xnor2_2 _0926_ (.A(_0286_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__xor2_4 _0927_ (.A(_0285_),
    .B(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__xnor2_4 _0928_ (.A(tdc_inst_capt_reg_r_1_2 ),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__xnor2_4 _0929_ (.A(_0281_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _0930_ (.A(tdc_inst_capt_reg_r_1_43 ),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0931_ (.A(tdc_inst_capt_reg_r_1_48 ),
    .Y(_0294_));
 sky130_fd_sc_hd__xor2_2 _0932_ (.A(tdc_inst_capt_reg_r_1_50 ),
    .B(tdc_inst_capt_reg_r_1_47 ),
    .X(_0295_));
 sky130_fd_sc_hd__xnor2_2 _0933_ (.A(tdc_inst_capt_reg_r_1_45 ),
    .B(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__xnor2_2 _0934_ (.A(_0294_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__xnor2_2 _0935_ (.A(_0293_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__or2_1 _0936_ (.A(tdc_inst_capt_reg_r_1_56 ),
    .B(tdc_inst_capt_reg_r_1_54 ),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _0937_ (.A(tdc_inst_capt_reg_r_1_56 ),
    .B(tdc_inst_capt_reg_r_1_54 ),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xor2_2 _0939_ (.A(tdc_inst_capt_reg_r_1_52 ),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(tdc_inst_capt_reg_r_1_1 ),
    .Y(_0303_));
 sky130_fd_sc_hd__xor2_2 _0941_ (.A(tdc_inst_capt_reg_r_1_62 ),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0304_));
 sky130_fd_sc_hd__xnor2_2 _0942_ (.A(tdc_inst_capt_reg_r_1_58 ),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__xnor2_2 _0943_ (.A(_0303_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__xor2_2 _0944_ (.A(_0302_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__xnor2_2 _0945_ (.A(tdc_inst_capt_reg_r_1_4 ),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__xor2_2 _0946_ (.A(_0298_),
    .B(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__xnor2_2 _0947_ (.A(tdc_inst_capt_reg_r_1_29 ),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__xor2_2 _0948_ (.A(_0292_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__xnor2_2 _0949_ (.A(tdc_inst_capt_reg_r_1_44 ),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__xor2_2 _0950_ (.A(_0280_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__xnor2_2 _0951_ (.A(tdc_inst_capt_reg_r_1_51 ),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__xor2_2 _0952_ (.A(_0253_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__xnor2_2 _0953_ (.A(tdc_inst_capt_reg_r_1_55 ),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_2 _0954_ (.A(_0222_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__xnor2_2 _0955_ (.A(_0221_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__xnor2_2 _0956_ (.A(_0220_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__nor2_1 _0957_ (.A(_0219_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__and2_1 _0958_ (.A(_0219_),
    .B(_0319_),
    .X(_0321_));
 sky130_fd_sc_hd__o21ai_1 _0959_ (.A1(_0320_),
    .A2(_0321_),
    .B1(_0218_),
    .Y(_0322_));
 sky130_fd_sc_hd__o211a_1 _0960_ (.A1(_0218_),
    .A2(uo_out[0]),
    .B1(_0073_),
    .C1(_0322_),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _0961_ (.A(tdc_inst_capt_reg_r_1_27 ),
    .B(_0234_),
    .X(_0323_));
 sky130_fd_sc_hd__a21o_1 _0962_ (.A1(tdc_inst_capt_reg_r_1_8 ),
    .A2(_0235_),
    .B1(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__o21ai_2 _0963_ (.A1(_0223_),
    .A2(_0252_),
    .B1(_0251_),
    .Y(_0325_));
 sky130_fd_sc_hd__or2_1 _0964_ (.A(_0237_),
    .B(_0247_),
    .X(_0326_));
 sky130_fd_sc_hd__o21a_1 _0965_ (.A1(_0236_),
    .A2(_0248_),
    .B1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__o21ai_2 _0966_ (.A1(_0254_),
    .A2(_0279_),
    .B1(_0278_),
    .Y(_0328_));
 sky130_fd_sc_hd__a21bo_1 _0967_ (.A1(tdc_inst_capt_reg_r_1_63 ),
    .A2(_0224_),
    .B1_N(_0225_),
    .X(_0329_));
 sky130_fd_sc_hd__a21bo_1 _0968_ (.A1(tdc_inst_capt_reg_r_1_41 ),
    .A2(_0229_),
    .B1_N(_0230_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _0969_ (.A(_0228_),
    .B(_0232_),
    .X(_0331_));
 sky130_fd_sc_hd__o21a_1 _0970_ (.A1(_0227_),
    .A2(_0233_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__xnor2_2 _0971_ (.A(_0330_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__xor2_2 _0972_ (.A(_0329_),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(_0241_),
    .B(_0243_),
    .X(_0335_));
 sky130_fd_sc_hd__o21ai_2 _0974_ (.A1(_0240_),
    .A2(_0244_),
    .B1(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__o21ai_2 _0975_ (.A1(_0261_),
    .A2(_0263_),
    .B1(_0266_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _0976_ (.A(tdc_inst_capt_reg_r_1_16 ),
    .B(tdc_inst_capt_reg_r_1_7 ),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _0977_ (.A(tdc_inst_capt_reg_r_1_22 ),
    .B(_0242_),
    .Y(_0339_));
 sky130_fd_sc_hd__a22oi_4 _0978_ (.A1(_0338_),
    .A2(_0339_),
    .B1(_0257_),
    .B2(_0259_),
    .Y(_0340_));
 sky130_fd_sc_hd__and4_1 _0979_ (.A(_0338_),
    .B(_0339_),
    .C(_0257_),
    .D(_0259_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _0980_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__xnor2_2 _0981_ (.A(_0337_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__xor2_2 _0982_ (.A(_0336_),
    .B(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _0983_ (.A(_0239_),
    .B(_0245_),
    .X(_0345_));
 sky130_fd_sc_hd__o21a_1 _0984_ (.A1(_0238_),
    .A2(_0246_),
    .B1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__xor2_2 _0985_ (.A(_0344_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__xnor2_2 _0986_ (.A(_0334_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_2 _0987_ (.A(_0328_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__xnor2_2 _0988_ (.A(_0327_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__or2_1 _0989_ (.A(_0268_),
    .B(_0274_),
    .X(_0351_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0275_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(_0267_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _0992_ (.A(tdc_inst_capt_reg_r_1_2 ),
    .B(_0290_),
    .Y(_0354_));
 sky130_fd_sc_hd__o21a_1 _0993_ (.A1(_0281_),
    .A2(_0291_),
    .B1(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _0994_ (.A(tdc_inst_capt_reg_r_1_15 ),
    .B(tdc_inst_capt_reg_r_1_0 ),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _0995_ (.A1(tdc_inst_capt_reg_r_1_11 ),
    .A2(_0262_),
    .B1(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__a21boi_1 _0996_ (.A1(tdc_inst_capt_reg_r_1_28 ),
    .A2(_0282_),
    .B1_N(_0283_),
    .Y(_0358_));
 sky130_fd_sc_hd__and2_1 _0997_ (.A(tdc_inst_capt_reg_r_1_26 ),
    .B(tdc_inst_capt_reg_r_1_23 ),
    .X(_0359_));
 sky130_fd_sc_hd__a21oi_1 _0998_ (.A1(tdc_inst_capt_reg_r_1_19 ),
    .A2(_0271_),
    .B1(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__or2_1 _0999_ (.A(_0358_),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _1000_ (.A(_0358_),
    .B(_0360_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0361_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__or2_1 _1002_ (.A(_0270_),
    .B(_0272_),
    .X(_0364_));
 sky130_fd_sc_hd__o21a_1 _1003_ (.A1(_0269_),
    .A2(_0273_),
    .B1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__xnor2_1 _1004_ (.A(_0363_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__xnor2_1 _1005_ (.A(_0357_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__xnor2_1 _1006_ (.A(_0355_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__and3_1 _1007_ (.A(_0351_),
    .B(_0353_),
    .C(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__a21o_1 _1008_ (.A1(_0351_),
    .A2(_0353_),
    .B1(_0368_),
    .X(_0370_));
 sky130_fd_sc_hd__and2b_1 _1009_ (.A_N(_0369_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(_0286_),
    .B(_0288_),
    .X(_0372_));
 sky130_fd_sc_hd__o21a_1 _1011_ (.A1(_0285_),
    .A2(_0289_),
    .B1(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(_0294_),
    .B(_0296_),
    .X(_0374_));
 sky130_fd_sc_hd__o21a_1 _1013_ (.A1(_0293_),
    .A2(_0297_),
    .B1(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _1014_ (.A(tdc_inst_capt_reg_r_1_42 ),
    .B(tdc_inst_capt_reg_r_1_38 ),
    .X(_0376_));
 sky130_fd_sc_hd__a21oi_2 _1015_ (.A1(tdc_inst_capt_reg_r_1_34 ),
    .A2(_0287_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__xor2_2 _1016_ (.A(_0375_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__xnor2_2 _1017_ (.A(_0373_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__a21boi_1 _1018_ (.A1(tdc_inst_capt_reg_r_1_52 ),
    .A2(_0299_),
    .B1_N(_0300_),
    .Y(_0380_));
 sky130_fd_sc_hd__and2_1 _1019_ (.A(tdc_inst_capt_reg_r_1_50 ),
    .B(tdc_inst_capt_reg_r_1_47 ),
    .X(_0381_));
 sky130_fd_sc_hd__a21oi_1 _1020_ (.A1(tdc_inst_capt_reg_r_1_45 ),
    .A2(_0295_),
    .B1(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__or2_1 _1021_ (.A(_0380_),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(_0380_),
    .B(_0382_),
    .Y(_0384_));
 sky130_fd_sc_hd__and2_1 _1023_ (.A(_0383_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _1024_ (.A(tdc_inst_capt_reg_r_1_62 ),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0386_));
 sky130_fd_sc_hd__a21o_1 _1025_ (.A1(tdc_inst_capt_reg_r_1_58 ),
    .A2(_0304_),
    .B1(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _1026_ (.A(_0303_),
    .B(_0305_),
    .X(_0388_));
 sky130_fd_sc_hd__o21a_1 _1027_ (.A1(_0302_),
    .A2(_0306_),
    .B1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__xnor2_2 _1028_ (.A(_0387_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__xnor2_2 _1029_ (.A(_0385_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _1030_ (.A(tdc_inst_capt_reg_r_1_4 ),
    .B(_0307_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21a_1 _1031_ (.A1(_0298_),
    .A2(_0308_),
    .B1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__xor2_2 _1032_ (.A(_0391_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__xnor2_2 _1033_ (.A(_0379_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(tdc_inst_capt_reg_r_1_29 ),
    .B(_0309_),
    .Y(_0396_));
 sky130_fd_sc_hd__o21ai_2 _1035_ (.A1(_0292_),
    .A2(_0310_),
    .B1(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__xnor2_2 _1036_ (.A(_0395_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__xnor2_2 _1037_ (.A(_0371_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _1038_ (.A(tdc_inst_capt_reg_r_1_44 ),
    .B(_0311_),
    .Y(_0400_));
 sky130_fd_sc_hd__o21ai_2 _1039_ (.A1(_0280_),
    .A2(_0312_),
    .B1(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_2 _1040_ (.A(_0399_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__xnor2_2 _1041_ (.A(_0350_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _1042_ (.A(tdc_inst_capt_reg_r_1_51 ),
    .B(_0313_),
    .Y(_0404_));
 sky130_fd_sc_hd__o21a_1 _1043_ (.A1(_0253_),
    .A2(_0314_),
    .B1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__xor2_2 _1044_ (.A(_0403_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__xnor2_2 _1045_ (.A(_0325_),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _1046_ (.A(tdc_inst_capt_reg_r_1_55 ),
    .B(_0315_),
    .Y(_0408_));
 sky130_fd_sc_hd__o21a_1 _1047_ (.A1(_0222_),
    .A2(_0316_),
    .B1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__xnor2_1 _1048_ (.A(_0407_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__xor2_1 _1049_ (.A(_0324_),
    .B(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _1050_ (.A(_0221_),
    .B(_0317_),
    .X(_0412_));
 sky130_fd_sc_hd__o21a_1 _1051_ (.A1(_0220_),
    .A2(_0318_),
    .B1(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__xor2_1 _1052_ (.A(_0411_),
    .B(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__xnor2_1 _1053_ (.A(_0320_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nand2_1 _1054_ (.A(_0218_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__o211a_1 _1055_ (.A1(_0218_),
    .A2(uo_out[1]),
    .B1(_0073_),
    .C1(_0416_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _1056_ (.A(_0407_),
    .B(_0409_),
    .X(_0417_));
 sky130_fd_sc_hd__or2b_1 _1057_ (.A(_0410_),
    .B_N(_0324_),
    .X(_0418_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0332_),
    .Y(_0419_));
 sky130_fd_sc_hd__and2_1 _1059_ (.A(_0329_),
    .B(_0333_),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_1 _1060_ (.A1(_0330_),
    .A2(_0419_),
    .B1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__or2b_1 _1061_ (.A(_0348_),
    .B_N(_0328_),
    .X(_0422_));
 sky130_fd_sc_hd__or2b_1 _1062_ (.A(_0327_),
    .B_N(_0349_),
    .X(_0423_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0422_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(_0344_),
    .B(_0346_),
    .Y(_0425_));
 sky130_fd_sc_hd__a21o_1 _1065_ (.A1(_0334_),
    .A2(_0347_),
    .B1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o21ai_1 _1066_ (.A1(_0355_),
    .A2(_0367_),
    .B1(_0370_),
    .Y(_0427_));
 sky130_fd_sc_hd__and2b_1 _1067_ (.A_N(_0343_),
    .B(_0336_),
    .X(_0428_));
 sky130_fd_sc_hd__a21oi_1 _1068_ (.A1(_0337_),
    .A2(_0342_),
    .B1(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__xnor2_1 _1069_ (.A(_0340_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__xor2_1 _1070_ (.A(_0427_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__xor2_1 _1071_ (.A(_0426_),
    .B(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__or2_1 _1072_ (.A(_0363_),
    .B(_0365_),
    .X(_0433_));
 sky130_fd_sc_hd__o21ai_1 _1073_ (.A1(_0357_),
    .A2(_0366_),
    .B1(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__and2b_1 _1074_ (.A_N(_0373_),
    .B(_0378_),
    .X(_0435_));
 sky130_fd_sc_hd__o21ba_1 _1075_ (.A1(_0375_),
    .A2(_0377_),
    .B1_N(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__xnor2_1 _1076_ (.A(_0361_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__xnor2_1 _1077_ (.A(_0434_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(_0387_),
    .Y(_0439_));
 sky130_fd_sc_hd__or2_1 _1079_ (.A(_0439_),
    .B(_0389_),
    .X(_0440_));
 sky130_fd_sc_hd__a21boi_1 _1080_ (.A1(_0385_),
    .A2(_0390_),
    .B1_N(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__nor2_1 _1081_ (.A(_0383_),
    .B(_0440_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_1 _1082_ (.A1(_0383_),
    .A2(_0441_),
    .B1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _1083_ (.A(_0391_),
    .B(_0393_),
    .Y(_0444_));
 sky130_fd_sc_hd__a21oi_1 _1084_ (.A1(_0379_),
    .A2(_0394_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__xnor2_1 _1085_ (.A(_0443_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__xnor2_1 _1086_ (.A(_0438_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__or2b_1 _1087_ (.A(_0395_),
    .B_N(_0397_),
    .X(_0448_));
 sky130_fd_sc_hd__a21boi_1 _1088_ (.A1(_0371_),
    .A2(_0398_),
    .B1_N(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__xor2_1 _1089_ (.A(_0447_),
    .B(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__xnor2_1 _1090_ (.A(_0432_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__and2b_1 _1091_ (.A_N(_0399_),
    .B(_0401_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1092_ (.A1(_0350_),
    .A2(_0402_),
    .B1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__xnor2_1 _1093_ (.A(_0451_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__xor2_1 _1094_ (.A(_0424_),
    .B(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _1095_ (.A(_0403_),
    .B(_0405_),
    .Y(_0456_));
 sky130_fd_sc_hd__a21oi_1 _1096_ (.A1(_0325_),
    .A2(_0406_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__xor2_1 _1097_ (.A(_0455_),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__xnor2_1 _1098_ (.A(_0421_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21oi_1 _1099_ (.A1(_0417_),
    .A2(_0418_),
    .B1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__and3_1 _1100_ (.A(_0417_),
    .B(_0418_),
    .C(_0459_),
    .X(_0461_));
 sky130_fd_sc_hd__nor2_1 _1101_ (.A(_0460_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nor2_1 _1102_ (.A(_0411_),
    .B(_0413_),
    .Y(_0463_));
 sky130_fd_sc_hd__a21o_1 _1103_ (.A1(_0320_),
    .A2(_0414_),
    .B1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__xnor2_1 _1104_ (.A(_0462_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _1105_ (.A(_0218_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__o211a_1 _1106_ (.A1(_0218_),
    .A2(uo_out[2]),
    .B1(_0073_),
    .C1(_0466_),
    .X(_0067_));
 sky130_fd_sc_hd__or2_1 _1107_ (.A(_0455_),
    .B(_0457_),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _1108_ (.A(_0421_),
    .B(_0458_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _1109_ (.A(_0427_),
    .B(_0430_),
    .Y(_0469_));
 sky130_fd_sc_hd__a21bo_1 _1110_ (.A1(_0426_),
    .A2(_0431_),
    .B1_N(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_1 _1111_ (.A(_0340_),
    .B(_0428_),
    .Y(_0471_));
 sky130_fd_sc_hd__or2b_1 _1112_ (.A(_0437_),
    .B_N(_0434_),
    .X(_0472_));
 sky130_fd_sc_hd__o21a_1 _1113_ (.A1(_0361_),
    .A2(_0436_),
    .B1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__or2_1 _1114_ (.A(_0471_),
    .B(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__nand2_1 _1115_ (.A(_0471_),
    .B(_0473_),
    .Y(_0475_));
 sky130_fd_sc_hd__and2_1 _1116_ (.A(_0474_),
    .B(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__and2_1 _1117_ (.A(_0438_),
    .B(_0446_),
    .X(_0477_));
 sky130_fd_sc_hd__nand2_1 _1118_ (.A(_0442_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__and2b_1 _1119_ (.A_N(_0445_),
    .B(_0443_),
    .X(_0479_));
 sky130_fd_sc_hd__or3_1 _1120_ (.A(_0442_),
    .B(_0479_),
    .C(_0477_),
    .X(_0480_));
 sky130_fd_sc_hd__and2_1 _1121_ (.A(_0478_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__xnor2_1 _1122_ (.A(_0476_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2_1 _1123_ (.A(_0447_),
    .B(_0449_),
    .Y(_0483_));
 sky130_fd_sc_hd__a21oi_1 _1124_ (.A1(_0432_),
    .A2(_0450_),
    .B1(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__xnor2_1 _1125_ (.A(_0482_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__xor2_1 _1126_ (.A(_0470_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__or2b_1 _1127_ (.A(_0454_),
    .B_N(_0424_),
    .X(_0487_));
 sky130_fd_sc_hd__o21a_1 _1128_ (.A1(_0451_),
    .A2(_0453_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__xnor2_1 _1129_ (.A(_0486_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__and3_1 _1130_ (.A(_0467_),
    .B(_0468_),
    .C(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__a21o_1 _1131_ (.A1(_0467_),
    .A2(_0468_),
    .B1(_0489_),
    .X(_0491_));
 sky130_fd_sc_hd__and2b_1 _1132_ (.A_N(_0490_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__a21oi_1 _1133_ (.A1(_0462_),
    .A2(_0464_),
    .B1(_0460_),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_1 _1134_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0075_),
    .Y(_0494_));
 sky130_fd_sc_hd__a21o_1 _1135_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__o211a_1 _1136_ (.A1(_0218_),
    .A2(uo_out[3]),
    .B1(_0073_),
    .C1(_0495_),
    .X(_0068_));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(_0486_),
    .B(_0488_),
    .X(_0496_));
 sky130_fd_sc_hd__and2b_1 _1138_ (.A_N(_0485_),
    .B(_0470_),
    .X(_0497_));
 sky130_fd_sc_hd__o21bai_1 _1139_ (.A1(_0482_),
    .A2(_0484_),
    .B1_N(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__a21bo_1 _1140_ (.A1(_0476_),
    .A2(_0480_),
    .B1_N(_0478_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1141_ (.A0(_0478_),
    .A1(_0499_),
    .S(_0474_),
    .X(_0500_));
 sky130_fd_sc_hd__xnor2_1 _1142_ (.A(_0498_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__and2_1 _1143_ (.A(_0496_),
    .B(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__nor2_1 _1144_ (.A(_0496_),
    .B(_0501_),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _1145_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__a21o_1 _1146_ (.A1(_0417_),
    .A2(_0418_),
    .B1(_0459_),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _1147_ (.A1(_0505_),
    .A2(_0491_),
    .B1(_0490_),
    .Y(_0506_));
 sky130_fd_sc_hd__a31o_1 _1148_ (.A1(_0462_),
    .A2(_0464_),
    .A3(_0492_),
    .B1(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__xnor2_1 _1149_ (.A(_0504_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(_0218_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__o211a_1 _1151_ (.A1(_0218_),
    .A2(uo_out[4]),
    .B1(_0073_),
    .C1(_0509_),
    .X(_0069_));
 sky130_fd_sc_hd__and2b_1 _1152_ (.A_N(_0075_),
    .B(uo_out[5]),
    .X(_0510_));
 sky130_fd_sc_hd__o2bb2a_1 _1153_ (.A1_N(_0498_),
    .A2_N(_0500_),
    .B1(_0474_),
    .B2(_0478_),
    .X(_0511_));
 sky130_fd_sc_hd__a21oi_1 _1154_ (.A1(_0504_),
    .A2(_0507_),
    .B1(_0503_),
    .Y(_0512_));
 sky130_fd_sc_hd__o21ai_1 _1155_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0075_),
    .Y(_0513_));
 sky130_fd_sc_hd__a21oi_1 _1156_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__o21a_1 _1157_ (.A1(_0510_),
    .A2(_0514_),
    .B1(_0073_),
    .X(_0070_));
 sky130_fd_sc_hd__o211a_1 _1158_ (.A1(uo_out[6]),
    .A2(_0218_),
    .B1(_0073_),
    .C1(_0513_),
    .X(_0071_));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(ui_in[0]),
    .D(_0000_),
    .Q(tdc_inst_pg_pg_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0001_),
    .Q(tdc_inst_capt_reg_r_1_0 ));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0002_),
    .Q(tdc_inst_capt_reg_r_1_1 ));
 sky130_fd_sc_hd__dfxtp_2 _1162_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0003_),
    .Q(tdc_inst_capt_reg_r_1_2 ));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0004_),
    .Q(tdc_inst_capt_reg_r_1_3 ));
 sky130_fd_sc_hd__dfxtp_2 _1164_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0005_),
    .Q(tdc_inst_capt_reg_r_1_4 ));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0006_),
    .Q(tdc_inst_capt_reg_r_1_5 ));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0007_),
    .Q(tdc_inst_capt_reg_r_1_6 ));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0008_),
    .Q(tdc_inst_capt_reg_r_1_7 ));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0009_),
    .Q(tdc_inst_capt_reg_r_1_8 ));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0010_),
    .Q(tdc_inst_capt_reg_r_1_9 ));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0011_),
    .Q(tdc_inst_capt_reg_r_1_10 ));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0012_),
    .Q(tdc_inst_capt_reg_r_1_11 ));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0013_),
    .Q(tdc_inst_capt_reg_r_1_12 ));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0014_),
    .Q(tdc_inst_capt_reg_r_1_13 ));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(_0015_),
    .Q(tdc_inst_capt_reg_r_1_14 ));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0016_),
    .Q(tdc_inst_capt_reg_r_1_15 ));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0017_),
    .Q(tdc_inst_capt_reg_r_1_16 ));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(_0018_),
    .Q(tdc_inst_capt_reg_r_1_17 ));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.CLK(clknet_4_10_0_ui_in[1]),
    .D(_0019_),
    .Q(tdc_inst_capt_reg_r_1_18 ));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(clknet_4_10_0_ui_in[1]),
    .D(_0020_),
    .Q(tdc_inst_capt_reg_r_1_19 ));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0021_),
    .Q(tdc_inst_capt_reg_r_1_20 ));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0022_),
    .Q(tdc_inst_capt_reg_r_1_21 ));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0023_),
    .Q(tdc_inst_capt_reg_r_1_22 ));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(clknet_4_8_0_ui_in[1]),
    .D(_0024_),
    .Q(tdc_inst_capt_reg_r_1_23 ));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0025_),
    .Q(tdc_inst_capt_reg_r_1_24 ));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0026_),
    .Q(tdc_inst_capt_reg_r_1_25 ));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.CLK(clknet_4_8_0_ui_in[1]),
    .D(_0027_),
    .Q(tdc_inst_capt_reg_r_1_26 ));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0028_),
    .Q(tdc_inst_capt_reg_r_1_27 ));
 sky130_fd_sc_hd__dfxtp_2 _1188_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0029_),
    .Q(tdc_inst_capt_reg_r_1_28 ));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0030_),
    .Q(tdc_inst_capt_reg_r_1_29 ));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(clknet_4_2_0_ui_in[1]),
    .D(_0031_),
    .Q(tdc_inst_capt_reg_r_1_30 ));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0032_),
    .Q(tdc_inst_capt_reg_r_1_31 ));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_4_2_0_ui_in[1]),
    .D(_0033_),
    .Q(tdc_inst_capt_reg_r_1_32 ));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0034_),
    .Q(tdc_inst_capt_reg_r_1_33 ));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.CLK(clknet_4_2_0_ui_in[1]),
    .D(_0035_),
    .Q(tdc_inst_capt_reg_r_1_34 ));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0036_),
    .Q(tdc_inst_capt_reg_r_1_35 ));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0037_),
    .Q(tdc_inst_capt_reg_r_1_36 ));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0038_),
    .Q(tdc_inst_capt_reg_r_1_37 ));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.CLK(clknet_4_2_0_ui_in[1]),
    .D(_0039_),
    .Q(tdc_inst_capt_reg_r_1_38 ));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0040_),
    .Q(tdc_inst_capt_reg_r_1_39 ));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0041_),
    .Q(tdc_inst_capt_reg_r_1_40 ));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0042_),
    .Q(tdc_inst_capt_reg_r_1_41 ));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(clknet_4_0_0_ui_in[1]),
    .D(_0043_),
    .Q(tdc_inst_capt_reg_r_1_42 ));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0044_),
    .Q(tdc_inst_capt_reg_r_1_43 ));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0045_),
    .Q(tdc_inst_capt_reg_r_1_44 ));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0046_),
    .Q(tdc_inst_capt_reg_r_1_45 ));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0047_),
    .Q(tdc_inst_capt_reg_r_1_46 ));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0048_),
    .Q(tdc_inst_capt_reg_r_1_47 ));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0049_),
    .Q(tdc_inst_capt_reg_r_1_48 ));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0050_),
    .Q(tdc_inst_capt_reg_r_1_49 ));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0051_),
    .Q(tdc_inst_capt_reg_r_1_50 ));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0052_),
    .Q(tdc_inst_capt_reg_r_1_51 ));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0053_),
    .Q(tdc_inst_capt_reg_r_1_52 ));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0054_),
    .Q(tdc_inst_capt_reg_r_1_53 ));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0055_),
    .Q(tdc_inst_capt_reg_r_1_54 ));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0056_),
    .Q(tdc_inst_capt_reg_r_1_55 ));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0057_),
    .Q(tdc_inst_capt_reg_r_1_56 ));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0058_),
    .Q(tdc_inst_capt_reg_r_1_57 ));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0059_),
    .Q(tdc_inst_capt_reg_r_1_58 ));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0060_),
    .Q(tdc_inst_capt_reg_r_1_59 ));
 sky130_fd_sc_hd__dfxtp_1 _1220_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0061_),
    .Q(tdc_inst_capt_reg_r_1_60 ));
 sky130_fd_sc_hd__dfxtp_1 _1221_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0062_),
    .Q(tdc_inst_capt_reg_r_1_61 ));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0063_),
    .Q(tdc_inst_capt_reg_r_1_62 ));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0064_),
    .Q(tdc_inst_capt_reg_r_1_63 ));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0065_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0066_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0067_),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0068_),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0069_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 _1229_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0070_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0071_),
    .Q(net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_ui_in_1  (.A(ui_in[1]),
    .X(clknet_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_0_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_10_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_11_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_12_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_13_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_14_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_15_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_1_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_2_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_3_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_4_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_5_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_6_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_7_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_8_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_9_0_ui_in[1]));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net1),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net16),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net16),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net16),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net11),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net11),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net11),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net177),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net186),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 hold11 (.A(net188),
    .X(uo_out[2]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net192),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 hold13 (.A(net194),
    .X(uo_out[3]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net183),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 hold15 (.A(net185),
    .X(uo_out[6]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net195),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 hold17 (.A(net178),
    .X(uo_out[5]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net197),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 hold19 (.A(net180),
    .X(uo_out[0]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net179),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net196),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 hold21 (.A(net182),
    .X(uo_out[1]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net165),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net175),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net176),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net167),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net171),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net172),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net166),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net169),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net181),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net170),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net168),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net173),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net174),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net198),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net199),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net200),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net162),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net164),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net163),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 hold4 (.A(net184),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 hold5 (.A(net190),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 hold6 (.A(net187),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 hold7 (.A(net193),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net189),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 hold9 (.A(net191),
    .X(uo_out[4]));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ena),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(ui_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_0_DFE  (.CLK(clknet_4_13_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_0 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_0 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_10_DFE  (.CLK(clknet_4_12_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_10 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_10 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_11_DFE  (.CLK(clknet_4_12_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_11 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_11 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_12_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_12 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_12 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_13_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_13 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_13 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_14_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_14 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_14 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_15_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_15 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_15 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_16_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_16 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_16 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_17_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_17 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_17 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_18_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_18 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_18 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_19_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_19 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_19 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_1_DFE  (.CLK(clknet_4_13_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_1 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_1 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_20_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_20 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_20 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_21_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_21 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_21 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_22_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_22 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_22 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_23_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_23 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_23 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_24_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_24 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_24 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_25_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_25 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_25 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_26_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_26 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_26 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_27_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_27 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_27 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_28_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_28 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_28 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_29_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_29 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_29 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_2_DFE  (.CLK(clknet_4_13_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_2 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_2 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_30_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_30 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_30 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_31_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_31 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_31 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_32_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_32 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_32 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_33_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_33 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_33 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_34_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_34 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_34 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_35_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_35 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_35 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_36_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_36 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_36 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_37_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_37 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_37 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_38_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_38 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_38 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_39_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_39 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_39 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_3_DFE  (.CLK(clknet_4_13_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_3 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_3 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_40_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_40 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_40 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_41_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_41 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_41 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_42_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_42 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_42 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_43_DFE  (.CLK(clknet_4_6_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_43 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_43 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_44_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_44 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_44 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_45_DFE  (.CLK(clknet_4_6_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_45 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_45 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_46_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_46 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_46 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_47_DFE  (.CLK(clknet_4_4_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_47 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_47 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_48_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_48 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_48 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_49_DFE  (.CLK(clknet_4_4_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_49 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_49 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_4_DFE  (.CLK(clknet_4_13_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_4 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_4 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_50_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_50 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_50 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_51_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_51 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_51 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_52_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_52 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_52 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_53_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_53 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_53 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_54_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_54 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_54 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_55_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_55 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_55 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_56_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_56 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_56 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_57_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_57 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_57 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_58_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_58 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_58 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_59_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_59 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_59 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_5_DFE  (.CLK(clknet_4_13_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_5 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_5 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_60_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_60 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_60 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_61_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_61 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_61 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_62_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_62 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_62 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_63_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_63 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_63 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_6_DFE  (.CLK(clknet_4_12_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_6 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_6 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_7_DFE  (.CLK(clknet_4_12_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_7 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_7 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_8_DFE  (.CLK(clknet_4_12_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_8 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_8 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_9_DFE  (.CLK(clknet_4_12_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_9 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_9 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_0_FA  (.A(net90),
    .B(net17),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_0 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_1 ),
    .SUM(tdc_inst_dl_capt_D_0 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_0_FA_17  (.LO(net17));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_0_FA_90  (.HI(net90));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_10_FA  (.A(net91),
    .B(net18),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_10 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_11 ),
    .SUM(tdc_inst_dl_capt_D_10 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_10_FA_18  (.LO(net18));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_10_FA_91  (.HI(net91));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_11_FA  (.A(net92),
    .B(net19),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_11 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_12 ),
    .SUM(tdc_inst_dl_capt_D_11 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_11_FA_19  (.LO(net19));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_11_FA_92  (.HI(net92));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_12_FA  (.A(net93),
    .B(net20),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_12 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_13 ),
    .SUM(tdc_inst_dl_capt_D_12 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_12_FA_20  (.LO(net20));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_12_FA_93  (.HI(net93));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_13_FA  (.A(net94),
    .B(net21),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_13 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_14 ),
    .SUM(tdc_inst_dl_capt_D_13 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_13_FA_21  (.LO(net21));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_13_FA_94  (.HI(net94));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_14_FA  (.A(net95),
    .B(net22),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_14 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_15 ),
    .SUM(tdc_inst_dl_capt_D_14 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_14_FA_22  (.LO(net22));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_14_FA_95  (.HI(net95));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_15_FA  (.A(net96),
    .B(net23),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_15 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_16 ),
    .SUM(tdc_inst_dl_capt_D_15 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_15_FA_23  (.LO(net23));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_15_FA_96  (.HI(net96));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_16_FA  (.A(net97),
    .B(net24),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_16 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_17 ),
    .SUM(tdc_inst_dl_capt_D_16 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_16_FA_24  (.LO(net24));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_16_FA_97  (.HI(net97));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_17_FA  (.A(net98),
    .B(net25),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_17 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_18 ),
    .SUM(tdc_inst_dl_capt_D_17 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_17_FA_25  (.LO(net25));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_17_FA_98  (.HI(net98));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_18_FA  (.A(net99),
    .B(net26),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_18 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_19 ),
    .SUM(tdc_inst_dl_capt_D_18 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_18_FA_26  (.LO(net26));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_18_FA_99  (.HI(net99));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_19_FA  (.A(net100),
    .B(net27),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_19 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_20 ),
    .SUM(tdc_inst_dl_capt_D_19 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_19_FA_100  (.HI(net100));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_19_FA_27  (.LO(net27));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_1_FA  (.A(net101),
    .B(net28),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_1 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_2 ),
    .SUM(tdc_inst_dl_capt_D_1 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_1_FA_101  (.HI(net101));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_1_FA_28  (.LO(net28));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_20_FA  (.A(net102),
    .B(net29),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_20 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_21 ),
    .SUM(tdc_inst_dl_capt_D_20 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_20_FA_102  (.HI(net102));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_20_FA_29  (.LO(net29));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_21_FA  (.A(net103),
    .B(net30),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_21 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_22 ),
    .SUM(tdc_inst_dl_capt_D_21 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_21_FA_103  (.HI(net103));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_21_FA_30  (.LO(net30));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_22_FA  (.A(net104),
    .B(net31),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_22 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_23 ),
    .SUM(tdc_inst_dl_capt_D_22 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_22_FA_104  (.HI(net104));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_22_FA_31  (.LO(net31));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_23_FA  (.A(net105),
    .B(net32),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_23 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_24 ),
    .SUM(tdc_inst_dl_capt_D_23 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_23_FA_105  (.HI(net105));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_23_FA_32  (.LO(net32));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_24_FA  (.A(net106),
    .B(net33),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_24 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_25 ),
    .SUM(tdc_inst_dl_capt_D_24 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_24_FA_106  (.HI(net106));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_24_FA_33  (.LO(net33));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_25_FA  (.A(net107),
    .B(net34),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_25 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_26 ),
    .SUM(tdc_inst_dl_capt_D_25 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_25_FA_107  (.HI(net107));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_25_FA_34  (.LO(net34));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_26_FA  (.A(net108),
    .B(net35),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_26 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_27 ),
    .SUM(tdc_inst_dl_capt_D_26 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_26_FA_108  (.HI(net108));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_26_FA_35  (.LO(net35));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_27_FA  (.A(net109),
    .B(net36),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_27 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_28 ),
    .SUM(tdc_inst_dl_capt_D_27 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_27_FA_109  (.HI(net109));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_27_FA_36  (.LO(net36));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_28_FA  (.A(net110),
    .B(net37),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_28 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_29 ),
    .SUM(tdc_inst_dl_capt_D_28 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_28_FA_110  (.HI(net110));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_28_FA_37  (.LO(net37));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_29_FA  (.A(net111),
    .B(net38),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_29 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_30 ),
    .SUM(tdc_inst_dl_capt_D_29 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_29_FA_111  (.HI(net111));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_29_FA_38  (.LO(net38));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_2_FA  (.A(net112),
    .B(net39),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_2 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_3 ),
    .SUM(tdc_inst_dl_capt_D_2 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_2_FA_112  (.HI(net112));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_2_FA_39  (.LO(net39));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_30_FA  (.A(net113),
    .B(net40),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_30 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_31 ),
    .SUM(tdc_inst_dl_capt_D_30 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_30_FA_113  (.HI(net113));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_30_FA_40  (.LO(net40));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_31_FA  (.A(net114),
    .B(net41),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_31 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_32 ),
    .SUM(tdc_inst_dl_capt_D_31 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_31_FA_114  (.HI(net114));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_31_FA_41  (.LO(net41));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_32_FA  (.A(net115),
    .B(net42),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_32 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_33 ),
    .SUM(tdc_inst_dl_capt_D_32 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_32_FA_115  (.HI(net115));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_32_FA_42  (.LO(net42));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_33_FA  (.A(net116),
    .B(net43),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_33 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_34 ),
    .SUM(tdc_inst_dl_capt_D_33 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_33_FA_116  (.HI(net116));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_33_FA_43  (.LO(net43));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_34_FA  (.A(net117),
    .B(net44),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_34 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_35 ),
    .SUM(tdc_inst_dl_capt_D_34 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_34_FA_117  (.HI(net117));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_34_FA_44  (.LO(net44));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_35_FA  (.A(net118),
    .B(net45),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_35 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_36 ),
    .SUM(tdc_inst_dl_capt_D_35 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_35_FA_118  (.HI(net118));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_35_FA_45  (.LO(net45));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_36_FA  (.A(net119),
    .B(net46),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_36 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_37 ),
    .SUM(tdc_inst_dl_capt_D_36 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_36_FA_119  (.HI(net119));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_36_FA_46  (.LO(net46));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_37_FA  (.A(net120),
    .B(net47),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_37 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_38 ),
    .SUM(tdc_inst_dl_capt_D_37 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_37_FA_120  (.HI(net120));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_37_FA_47  (.LO(net47));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_38_FA  (.A(net121),
    .B(net48),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_38 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_39 ),
    .SUM(tdc_inst_dl_capt_D_38 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_38_FA_121  (.HI(net121));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_38_FA_48  (.LO(net48));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_39_FA  (.A(net122),
    .B(net49),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_39 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_40 ),
    .SUM(tdc_inst_dl_capt_D_39 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_39_FA_122  (.HI(net122));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_39_FA_49  (.LO(net49));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_3_FA  (.A(net123),
    .B(net50),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_3 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_4 ),
    .SUM(tdc_inst_dl_capt_D_3 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_3_FA_123  (.HI(net123));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_3_FA_50  (.LO(net50));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_40_FA  (.A(net124),
    .B(net51),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_40 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_41 ),
    .SUM(tdc_inst_dl_capt_D_40 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_40_FA_124  (.HI(net124));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_40_FA_51  (.LO(net51));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_41_FA  (.A(net125),
    .B(net52),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_41 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_42 ),
    .SUM(tdc_inst_dl_capt_D_41 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_41_FA_125  (.HI(net125));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_41_FA_52  (.LO(net52));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_42_FA  (.A(net126),
    .B(net53),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_42 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_43 ),
    .SUM(tdc_inst_dl_capt_D_42 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_42_FA_126  (.HI(net126));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_42_FA_53  (.LO(net53));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_43_FA  (.A(net127),
    .B(net54),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_43 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_44 ),
    .SUM(tdc_inst_dl_capt_D_43 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_43_FA_127  (.HI(net127));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_43_FA_54  (.LO(net54));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_44_FA  (.A(net128),
    .B(net55),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_44 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_45 ),
    .SUM(tdc_inst_dl_capt_D_44 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_44_FA_128  (.HI(net128));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_44_FA_55  (.LO(net55));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_45_FA  (.A(net129),
    .B(net56),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_45 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_46 ),
    .SUM(tdc_inst_dl_capt_D_45 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_45_FA_129  (.HI(net129));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_45_FA_56  (.LO(net56));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_46_FA  (.A(net130),
    .B(net57),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_46 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_47 ),
    .SUM(tdc_inst_dl_capt_D_46 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_46_FA_130  (.HI(net130));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_46_FA_57  (.LO(net57));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_47_FA  (.A(net131),
    .B(net58),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_47 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_48 ),
    .SUM(tdc_inst_dl_capt_D_47 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_47_FA_131  (.HI(net131));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_47_FA_58  (.LO(net58));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_48_FA  (.A(net132),
    .B(net59),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_48 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_49 ),
    .SUM(tdc_inst_dl_capt_D_48 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_48_FA_132  (.HI(net132));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_48_FA_59  (.LO(net59));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_49_FA  (.A(net133),
    .B(net60),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_49 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_50 ),
    .SUM(tdc_inst_dl_capt_D_49 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_49_FA_133  (.HI(net133));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_49_FA_60  (.LO(net60));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_4_FA  (.A(net134),
    .B(net61),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_4 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_5 ),
    .SUM(tdc_inst_dl_capt_D_4 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_4_FA_134  (.HI(net134));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_4_FA_61  (.LO(net61));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_50_FA  (.A(net135),
    .B(net62),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_50 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_51 ),
    .SUM(tdc_inst_dl_capt_D_50 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_50_FA_135  (.HI(net135));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_50_FA_62  (.LO(net62));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_51_FA  (.A(net136),
    .B(net63),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_51 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_52 ),
    .SUM(tdc_inst_dl_capt_D_51 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_51_FA_136  (.HI(net136));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_51_FA_63  (.LO(net63));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_52_FA  (.A(net137),
    .B(net64),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_52 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_53 ),
    .SUM(tdc_inst_dl_capt_D_52 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_52_FA_137  (.HI(net137));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_52_FA_64  (.LO(net64));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_53_FA  (.A(net138),
    .B(net65),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_53 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_54 ),
    .SUM(tdc_inst_dl_capt_D_53 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_53_FA_138  (.HI(net138));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_53_FA_65  (.LO(net65));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_54_FA  (.A(net139),
    .B(net66),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_54 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_55 ),
    .SUM(tdc_inst_dl_capt_D_54 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_54_FA_139  (.HI(net139));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_54_FA_66  (.LO(net66));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_55_FA  (.A(net140),
    .B(net67),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_55 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_56 ),
    .SUM(tdc_inst_dl_capt_D_55 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_55_FA_140  (.HI(net140));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_55_FA_67  (.LO(net67));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_56_FA  (.A(net141),
    .B(net68),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_56 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_57 ),
    .SUM(tdc_inst_dl_capt_D_56 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_56_FA_141  (.HI(net141));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_56_FA_68  (.LO(net68));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_57_FA  (.A(net142),
    .B(net69),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_57 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_58 ),
    .SUM(tdc_inst_dl_capt_D_57 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_57_FA_142  (.HI(net142));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_57_FA_69  (.LO(net69));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_58_FA  (.A(net143),
    .B(net70),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_58 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_59 ),
    .SUM(tdc_inst_dl_capt_D_58 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_58_FA_143  (.HI(net143));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_58_FA_70  (.LO(net70));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_59_FA  (.A(net144),
    .B(net71),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_59 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_60 ),
    .SUM(tdc_inst_dl_capt_D_59 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_59_FA_144  (.HI(net144));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_59_FA_71  (.LO(net71));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_5_FA  (.A(net145),
    .B(net72),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_5 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_6 ),
    .SUM(tdc_inst_dl_capt_D_5 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_5_FA_145  (.HI(net145));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_5_FA_72  (.LO(net72));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_60_FA  (.A(net146),
    .B(net73),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_60 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_61 ),
    .SUM(tdc_inst_dl_capt_D_60 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_60_FA_146  (.HI(net146));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_60_FA_73  (.LO(net73));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_61_FA  (.A(net147),
    .B(net74),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_61 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_62 ),
    .SUM(tdc_inst_dl_capt_D_61 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_61_FA_147  (.HI(net147));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_61_FA_74  (.LO(net74));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_62_FA  (.A(net148),
    .B(net75),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_62 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_63 ),
    .SUM(tdc_inst_dl_capt_D_62 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_62_FA_148  (.HI(net148));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_62_FA_75  (.LO(net75));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_63_FA  (.A(net149),
    .B(net76),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_63 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_keep_co ),
    .SUM(tdc_inst_dl_capt_D_63 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_63_FA_149  (.HI(net149));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_63_FA_76  (.LO(net76));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_6_FA  (.A(net150),
    .B(net77),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_6 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_7 ),
    .SUM(tdc_inst_dl_capt_D_6 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_6_FA_150  (.HI(net150));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_6_FA_77  (.LO(net77));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_7_FA  (.A(net151),
    .B(net78),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_7 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_8 ),
    .SUM(tdc_inst_dl_capt_D_7 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_7_FA_151  (.HI(net151));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_7_FA_78  (.LO(net78));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_8_FA  (.A(net152),
    .B(net79),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_8 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_9 ),
    .SUM(tdc_inst_dl_capt_D_8 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_8_FA_152  (.HI(net152));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_8_FA_79  (.LO(net79));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_9_FA  (.A(net153),
    .B(net80),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_9 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_10 ),
    .SUM(tdc_inst_dl_capt_D_9 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_9_FA_153  (.HI(net153));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_9_FA_80  (.LO(net80));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_154 (.HI(net154));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_155 (.HI(net155));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_156 (.HI(net156));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_157 (.HI(net157));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_158 (.HI(net158));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_159 (.HI(net159));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_160 (.HI(net160));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_161 (.HI(net161));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_89 (.LO(net89));
 assign uio_oe[0] = net154;
 assign uio_oe[1] = net155;
 assign uio_oe[2] = net156;
 assign uio_oe[3] = net157;
 assign uio_oe[4] = net158;
 assign uio_oe[5] = net159;
 assign uio_oe[6] = net160;
 assign uio_oe[7] = net161;
 assign uio_out[0] = net81;
 assign uio_out[1] = net82;
 assign uio_out[2] = net83;
 assign uio_out[3] = net84;
 assign uio_out[4] = net85;
 assign uio_out[5] = net86;
 assign uio_out[6] = net87;
 assign uio_out[7] = net88;
 assign uo_out[7] = net89;
endmodule

