// This is the unpowered netlist.
module tt_um_hsc_tdc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net2;
 wire net3;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire tdc_inst_capt_out_0 ;
 wire tdc_inst_capt_out_10 ;
 wire tdc_inst_capt_out_11 ;
 wire tdc_inst_capt_out_12 ;
 wire tdc_inst_capt_out_13 ;
 wire tdc_inst_capt_out_14 ;
 wire tdc_inst_capt_out_15 ;
 wire tdc_inst_capt_out_16 ;
 wire tdc_inst_capt_out_17 ;
 wire tdc_inst_capt_out_18 ;
 wire tdc_inst_capt_out_19 ;
 wire tdc_inst_capt_out_1 ;
 wire tdc_inst_capt_out_20 ;
 wire tdc_inst_capt_out_21 ;
 wire tdc_inst_capt_out_22 ;
 wire tdc_inst_capt_out_23 ;
 wire tdc_inst_capt_out_24 ;
 wire tdc_inst_capt_out_25 ;
 wire tdc_inst_capt_out_26 ;
 wire tdc_inst_capt_out_27 ;
 wire tdc_inst_capt_out_28 ;
 wire tdc_inst_capt_out_29 ;
 wire tdc_inst_capt_out_2 ;
 wire tdc_inst_capt_out_30 ;
 wire tdc_inst_capt_out_31 ;
 wire tdc_inst_capt_out_32 ;
 wire tdc_inst_capt_out_33 ;
 wire tdc_inst_capt_out_34 ;
 wire tdc_inst_capt_out_35 ;
 wire tdc_inst_capt_out_36 ;
 wire tdc_inst_capt_out_37 ;
 wire tdc_inst_capt_out_38 ;
 wire tdc_inst_capt_out_39 ;
 wire tdc_inst_capt_out_3 ;
 wire tdc_inst_capt_out_40 ;
 wire tdc_inst_capt_out_41 ;
 wire tdc_inst_capt_out_42 ;
 wire tdc_inst_capt_out_43 ;
 wire tdc_inst_capt_out_44 ;
 wire tdc_inst_capt_out_45 ;
 wire tdc_inst_capt_out_46 ;
 wire tdc_inst_capt_out_47 ;
 wire tdc_inst_capt_out_48 ;
 wire tdc_inst_capt_out_49 ;
 wire tdc_inst_capt_out_4 ;
 wire tdc_inst_capt_out_50 ;
 wire tdc_inst_capt_out_51 ;
 wire tdc_inst_capt_out_52 ;
 wire tdc_inst_capt_out_53 ;
 wire tdc_inst_capt_out_54 ;
 wire tdc_inst_capt_out_55 ;
 wire tdc_inst_capt_out_56 ;
 wire tdc_inst_capt_out_57 ;
 wire tdc_inst_capt_out_58 ;
 wire tdc_inst_capt_out_59 ;
 wire tdc_inst_capt_out_5 ;
 wire tdc_inst_capt_out_60 ;
 wire tdc_inst_capt_out_61 ;
 wire tdc_inst_capt_out_62 ;
 wire tdc_inst_capt_out_63 ;
 wire tdc_inst_capt_out_6 ;
 wire tdc_inst_capt_out_7 ;
 wire tdc_inst_capt_out_8 ;
 wire tdc_inst_capt_out_9 ;
 wire tdc_inst_capt_reg_r_1_0 ;
 wire tdc_inst_capt_reg_r_1_10 ;
 wire tdc_inst_capt_reg_r_1_11 ;
 wire tdc_inst_capt_reg_r_1_12 ;
 wire tdc_inst_capt_reg_r_1_13 ;
 wire tdc_inst_capt_reg_r_1_14 ;
 wire tdc_inst_capt_reg_r_1_15 ;
 wire tdc_inst_capt_reg_r_1_16 ;
 wire tdc_inst_capt_reg_r_1_17 ;
 wire tdc_inst_capt_reg_r_1_18 ;
 wire tdc_inst_capt_reg_r_1_19 ;
 wire tdc_inst_capt_reg_r_1_1 ;
 wire tdc_inst_capt_reg_r_1_20 ;
 wire tdc_inst_capt_reg_r_1_21 ;
 wire tdc_inst_capt_reg_r_1_22 ;
 wire tdc_inst_capt_reg_r_1_23 ;
 wire tdc_inst_capt_reg_r_1_24 ;
 wire tdc_inst_capt_reg_r_1_25 ;
 wire tdc_inst_capt_reg_r_1_26 ;
 wire tdc_inst_capt_reg_r_1_27 ;
 wire tdc_inst_capt_reg_r_1_28 ;
 wire tdc_inst_capt_reg_r_1_29 ;
 wire tdc_inst_capt_reg_r_1_2 ;
 wire tdc_inst_capt_reg_r_1_30 ;
 wire tdc_inst_capt_reg_r_1_31 ;
 wire tdc_inst_capt_reg_r_1_32 ;
 wire tdc_inst_capt_reg_r_1_33 ;
 wire tdc_inst_capt_reg_r_1_34 ;
 wire tdc_inst_capt_reg_r_1_35 ;
 wire tdc_inst_capt_reg_r_1_36 ;
 wire tdc_inst_capt_reg_r_1_37 ;
 wire tdc_inst_capt_reg_r_1_38 ;
 wire tdc_inst_capt_reg_r_1_39 ;
 wire tdc_inst_capt_reg_r_1_3 ;
 wire tdc_inst_capt_reg_r_1_40 ;
 wire tdc_inst_capt_reg_r_1_41 ;
 wire tdc_inst_capt_reg_r_1_42 ;
 wire tdc_inst_capt_reg_r_1_43 ;
 wire tdc_inst_capt_reg_r_1_44 ;
 wire tdc_inst_capt_reg_r_1_45 ;
 wire tdc_inst_capt_reg_r_1_46 ;
 wire tdc_inst_capt_reg_r_1_47 ;
 wire tdc_inst_capt_reg_r_1_48 ;
 wire tdc_inst_capt_reg_r_1_49 ;
 wire tdc_inst_capt_reg_r_1_4 ;
 wire tdc_inst_capt_reg_r_1_50 ;
 wire tdc_inst_capt_reg_r_1_51 ;
 wire tdc_inst_capt_reg_r_1_52 ;
 wire tdc_inst_capt_reg_r_1_53 ;
 wire tdc_inst_capt_reg_r_1_54 ;
 wire tdc_inst_capt_reg_r_1_55 ;
 wire tdc_inst_capt_reg_r_1_56 ;
 wire tdc_inst_capt_reg_r_1_57 ;
 wire tdc_inst_capt_reg_r_1_58 ;
 wire tdc_inst_capt_reg_r_1_59 ;
 wire tdc_inst_capt_reg_r_1_5 ;
 wire tdc_inst_capt_reg_r_1_60 ;
 wire tdc_inst_capt_reg_r_1_61 ;
 wire tdc_inst_capt_reg_r_1_62 ;
 wire tdc_inst_capt_reg_r_1_63 ;
 wire tdc_inst_capt_reg_r_1_6 ;
 wire tdc_inst_capt_reg_r_1_7 ;
 wire tdc_inst_capt_reg_r_1_8 ;
 wire tdc_inst_capt_reg_r_1_9 ;
 wire tdc_inst_dl_capt_D_0 ;
 wire tdc_inst_dl_capt_D_10 ;
 wire tdc_inst_dl_capt_D_11 ;
 wire tdc_inst_dl_capt_D_12 ;
 wire tdc_inst_dl_capt_D_13 ;
 wire tdc_inst_dl_capt_D_14 ;
 wire tdc_inst_dl_capt_D_15 ;
 wire tdc_inst_dl_capt_D_16 ;
 wire tdc_inst_dl_capt_D_17 ;
 wire tdc_inst_dl_capt_D_18 ;
 wire tdc_inst_dl_capt_D_19 ;
 wire tdc_inst_dl_capt_D_1 ;
 wire tdc_inst_dl_capt_D_20 ;
 wire tdc_inst_dl_capt_D_21 ;
 wire tdc_inst_dl_capt_D_22 ;
 wire tdc_inst_dl_capt_D_23 ;
 wire tdc_inst_dl_capt_D_24 ;
 wire tdc_inst_dl_capt_D_25 ;
 wire tdc_inst_dl_capt_D_26 ;
 wire tdc_inst_dl_capt_D_27 ;
 wire tdc_inst_dl_capt_D_28 ;
 wire tdc_inst_dl_capt_D_29 ;
 wire tdc_inst_dl_capt_D_2 ;
 wire tdc_inst_dl_capt_D_30 ;
 wire tdc_inst_dl_capt_D_31 ;
 wire tdc_inst_dl_capt_D_32 ;
 wire tdc_inst_dl_capt_D_33 ;
 wire tdc_inst_dl_capt_D_34 ;
 wire tdc_inst_dl_capt_D_35 ;
 wire tdc_inst_dl_capt_D_36 ;
 wire tdc_inst_dl_capt_D_37 ;
 wire tdc_inst_dl_capt_D_38 ;
 wire tdc_inst_dl_capt_D_39 ;
 wire tdc_inst_dl_capt_D_3 ;
 wire tdc_inst_dl_capt_D_40 ;
 wire tdc_inst_dl_capt_D_41 ;
 wire tdc_inst_dl_capt_D_42 ;
 wire tdc_inst_dl_capt_D_43 ;
 wire tdc_inst_dl_capt_D_44 ;
 wire tdc_inst_dl_capt_D_45 ;
 wire tdc_inst_dl_capt_D_46 ;
 wire tdc_inst_dl_capt_D_47 ;
 wire tdc_inst_dl_capt_D_48 ;
 wire tdc_inst_dl_capt_D_49 ;
 wire tdc_inst_dl_capt_D_4 ;
 wire tdc_inst_dl_capt_D_50 ;
 wire tdc_inst_dl_capt_D_51 ;
 wire tdc_inst_dl_capt_D_52 ;
 wire tdc_inst_dl_capt_D_53 ;
 wire tdc_inst_dl_capt_D_54 ;
 wire tdc_inst_dl_capt_D_55 ;
 wire tdc_inst_dl_capt_D_56 ;
 wire tdc_inst_dl_capt_D_57 ;
 wire tdc_inst_dl_capt_D_58 ;
 wire tdc_inst_dl_capt_D_59 ;
 wire tdc_inst_dl_capt_D_5 ;
 wire tdc_inst_dl_capt_D_60 ;
 wire tdc_inst_dl_capt_D_61 ;
 wire tdc_inst_dl_capt_D_62 ;
 wire tdc_inst_dl_capt_D_63 ;
 wire tdc_inst_dl_capt_D_6 ;
 wire tdc_inst_dl_capt_D_7 ;
 wire tdc_inst_dl_capt_D_8 ;
 wire tdc_inst_dl_capt_D_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_0 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_10 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_11 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_12 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_13 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_14 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_15 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_16 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_17 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_18 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_19 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_1 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_20 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_21 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_22 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_23 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_24 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_25 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_26 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_27 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_28 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_29 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_2 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_30 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_31 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_32 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_33 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_34 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_35 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_36 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_37 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_38 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_39 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_3 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_40 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_41 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_42 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_43 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_44 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_45 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_46 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_47 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_48 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_49 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_4 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_50 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_51 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_52 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_53 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_54 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_55 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_56 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_57 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_58 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_59 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_5 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_60 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_61 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_62 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_63 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_6 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_7 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_8 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_0 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_10 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_11 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_12 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_13 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_14 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_15 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_16 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_17 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_18 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_19 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_1 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_20 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_21 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_22 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_23 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_24 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_25 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_26 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_27 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_28 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_29 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_2 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_30 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_31 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_32 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_33 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_34 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_35 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_36 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_37 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_38 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_39 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_3 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_40 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_41 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_42 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_43 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_44 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_45 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_46 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_47 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_48 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_49 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_4 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_50 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_51 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_52 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_53 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_54 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_55 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_56 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_57 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_58 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_59 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_5 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_60 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_61 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_62 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_63 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_6 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_7 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_8 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_b_int_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_0 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_10 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_11 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_12 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_13 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_14 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_15 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_16 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_17 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_18 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_19 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_1 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_20 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_21 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_22 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_23 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_24 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_25 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_26 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_27 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_28 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_29 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_2 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_30 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_31 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_32 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_33 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_34 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_35 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_36 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_37 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_38 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_39 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_3 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_40 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_41 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_42 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_43 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_44 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_45 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_46 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_47 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_48 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_49 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_4 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_50 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_51 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_52 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_53 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_54 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_55 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_56 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_57 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_58 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_59 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_5 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_60 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_61 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_62 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_63 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_64 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_6 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_7 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_8 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_c_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_co ;
 wire tdc_inst_pc_inst_val_in ;
 wire tdc_inst_pc_inst_val_out ;
 wire tdc_inst_pg_pg_r_out ;
 wire tdc_inst_pg_val_r_out ;
 wire tdc_inst_pg_out ;
 wire tdc_inst_val_out_capt ;
 wire [1:0] clknet_0_ui_in;
 wire [0:0] clknet_1_0__leaf_ui_in;
 wire [0:0] clknet_1_1__leaf_ui_in;
 wire [1:0] clknet_4_0_0_ui_in;
 wire [1:0] clknet_4_10_0_ui_in;
 wire [1:0] clknet_4_11_0_ui_in;
 wire [1:0] clknet_4_12_0_ui_in;
 wire [1:0] clknet_4_13_0_ui_in;
 wire [1:0] clknet_4_14_0_ui_in;
 wire [1:0] clknet_4_15_0_ui_in;
 wire [1:0] clknet_4_1_0_ui_in;
 wire [1:0] clknet_4_2_0_ui_in;
 wire [1:0] clknet_4_3_0_ui_in;
 wire [1:0] clknet_4_4_0_ui_in;
 wire [1:0] clknet_4_5_0_ui_in;
 wire [1:0] clknet_4_6_0_ui_in;
 wire [1:0] clknet_4_7_0_ui_in;
 wire [1:0] clknet_4_8_0_ui_in;
 wire [1:0] clknet_4_9_0_ui_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net2));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__mux2_1 _0529_ (.A0(tdc_inst_pg_pg_r_out ),
    .A1(net6),
    .S(net4),
    .X(_0076_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0530_ (.A(_0076_),
    .X(tdc_inst_dl_inst_dl_genblk_dl_c_0 ));
 sky130_fd_sc_hd__clkbuf_4 _0531_ (.A(net2),
    .X(_0077_));
 sky130_fd_sc_hd__buf_2 _0532_ (.A(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0533_ (.A0(net5),
    .A1(net6),
    .S(net3),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_4 _0534_ (.A(net8),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_4 _0535_ (.A(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0536_ (.A0(tdc_inst_pg_pg_r_out ),
    .A1(_0079_),
    .S(_0081_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _0537_ (.A(_0078_),
    .B(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_1 _0538_ (.A(_0083_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _0539_ (.A0(tdc_inst_pg_val_r_out ),
    .A1(net7),
    .S(_0081_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _0540_ (.A(_0078_),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0541_ (.A(_0085_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0542_ (.A0(net33),
    .A1(net7),
    .S(net4),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0543_ (.A0(tdc_inst_val_out_capt ),
    .A1(_0086_),
    .S(_0081_),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _0544_ (.A(_0078_),
    .B(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0545_ (.A(_0088_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_2 _0546_ (.A(_0077_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0547_ (.A0(tdc_inst_capt_reg_r_1_0 ),
    .A1(tdc_inst_capt_out_0 ),
    .S(_0081_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _0548_ (.A(_0089_),
    .B(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _0549_ (.A(_0091_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0550_ (.A0(tdc_inst_capt_reg_r_1_1 ),
    .A1(tdc_inst_capt_out_1 ),
    .S(_0081_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _0551_ (.A(_0089_),
    .B(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_1 _0552_ (.A(_0093_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0553_ (.A0(tdc_inst_capt_reg_r_1_2 ),
    .A1(tdc_inst_capt_out_2 ),
    .S(_0081_),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _0554_ (.A(_0089_),
    .B(_0094_),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _0555_ (.A(_0095_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_4 _0556_ (.A(_0080_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0557_ (.A0(tdc_inst_capt_reg_r_1_3 ),
    .A1(tdc_inst_capt_out_3 ),
    .S(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _0558_ (.A(_0089_),
    .B(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0559_ (.A(_0098_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0560_ (.A0(tdc_inst_capt_reg_r_1_4 ),
    .A1(tdc_inst_capt_out_4 ),
    .S(_0096_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _0561_ (.A(_0089_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0562_ (.A(_0100_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0563_ (.A0(tdc_inst_capt_reg_r_1_5 ),
    .A1(tdc_inst_capt_out_5 ),
    .S(_0096_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _0564_ (.A(_0089_),
    .B(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _0565_ (.A(_0102_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0566_ (.A0(tdc_inst_capt_reg_r_1_6 ),
    .A1(tdc_inst_capt_out_6 ),
    .S(_0096_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _0567_ (.A(_0089_),
    .B(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0568_ (.A(_0104_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0569_ (.A0(tdc_inst_capt_reg_r_1_7 ),
    .A1(tdc_inst_capt_out_7 ),
    .S(_0096_),
    .X(_0105_));
 sky130_fd_sc_hd__and2_1 _0570_ (.A(_0089_),
    .B(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0571_ (.A(_0106_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0572_ (.A0(tdc_inst_capt_reg_r_1_8 ),
    .A1(tdc_inst_capt_out_8 ),
    .S(_0096_),
    .X(_0107_));
 sky130_fd_sc_hd__and2_1 _0573_ (.A(_0089_),
    .B(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0574_ (.A(_0108_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0575_ (.A0(tdc_inst_capt_reg_r_1_9 ),
    .A1(tdc_inst_capt_out_9 ),
    .S(_0096_),
    .X(_0109_));
 sky130_fd_sc_hd__and2_1 _0576_ (.A(_0089_),
    .B(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0577_ (.A(_0110_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_2 _0578_ (.A(_0077_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(tdc_inst_capt_reg_r_1_10 ),
    .A1(tdc_inst_capt_out_10 ),
    .S(_0096_),
    .X(_0112_));
 sky130_fd_sc_hd__and2_1 _0580_ (.A(_0111_),
    .B(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _0581_ (.A(_0113_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0582_ (.A0(tdc_inst_capt_reg_r_1_11 ),
    .A1(tdc_inst_capt_out_11 ),
    .S(_0096_),
    .X(_0114_));
 sky130_fd_sc_hd__and2_1 _0583_ (.A(_0111_),
    .B(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_1 _0584_ (.A(_0115_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(tdc_inst_capt_reg_r_1_12 ),
    .A1(tdc_inst_capt_out_12 ),
    .S(_0096_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _0586_ (.A(_0111_),
    .B(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _0587_ (.A(_0117_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _0588_ (.A(_0080_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(tdc_inst_capt_reg_r_1_13 ),
    .A1(tdc_inst_capt_out_13 ),
    .S(_0118_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _0590_ (.A(_0111_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0591_ (.A(_0120_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(tdc_inst_capt_reg_r_1_14 ),
    .A1(tdc_inst_capt_out_14 ),
    .S(_0118_),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _0593_ (.A(_0111_),
    .B(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _0594_ (.A(_0122_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(tdc_inst_capt_reg_r_1_15 ),
    .A1(tdc_inst_capt_out_15 ),
    .S(_0118_),
    .X(_0123_));
 sky130_fd_sc_hd__and2_1 _0596_ (.A(_0111_),
    .B(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0124_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(tdc_inst_capt_reg_r_1_16 ),
    .A1(tdc_inst_capt_out_16 ),
    .S(_0118_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _0599_ (.A(_0111_),
    .B(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0600_ (.A(_0126_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(tdc_inst_capt_reg_r_1_17 ),
    .A1(tdc_inst_capt_out_17 ),
    .S(_0118_),
    .X(_0127_));
 sky130_fd_sc_hd__and2_1 _0602_ (.A(_0111_),
    .B(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _0603_ (.A(_0128_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(tdc_inst_capt_reg_r_1_18 ),
    .A1(tdc_inst_capt_out_18 ),
    .S(_0118_),
    .X(_0129_));
 sky130_fd_sc_hd__and2_1 _0605_ (.A(_0111_),
    .B(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_1 _0606_ (.A(_0130_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0607_ (.A0(tdc_inst_capt_reg_r_1_19 ),
    .A1(tdc_inst_capt_out_19 ),
    .S(_0118_),
    .X(_0131_));
 sky130_fd_sc_hd__and2_1 _0608_ (.A(_0111_),
    .B(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0609_ (.A(_0132_),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_2 _0610_ (.A(_0077_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0611_ (.A0(tdc_inst_capt_reg_r_1_20 ),
    .A1(tdc_inst_capt_out_20 ),
    .S(_0118_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _0612_ (.A(_0133_),
    .B(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _0613_ (.A(_0135_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(tdc_inst_capt_reg_r_1_21 ),
    .A1(tdc_inst_capt_out_21 ),
    .S(_0118_),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _0615_ (.A(_0133_),
    .B(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0137_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0617_ (.A0(tdc_inst_capt_reg_r_1_22 ),
    .A1(tdc_inst_capt_out_22 ),
    .S(_0118_),
    .X(_0138_));
 sky130_fd_sc_hd__and2_1 _0618_ (.A(_0133_),
    .B(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _0619_ (.A(_0139_),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_4 _0620_ (.A(_0080_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0621_ (.A0(tdc_inst_capt_reg_r_1_23 ),
    .A1(tdc_inst_capt_out_23 ),
    .S(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _0622_ (.A(_0133_),
    .B(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0623_ (.A(_0142_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(tdc_inst_capt_reg_r_1_24 ),
    .A1(tdc_inst_capt_out_24 ),
    .S(_0140_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(_0133_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0626_ (.A(_0144_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(tdc_inst_capt_reg_r_1_25 ),
    .A1(tdc_inst_capt_out_25 ),
    .S(_0140_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _0628_ (.A(_0133_),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0629_ (.A(_0146_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(tdc_inst_capt_reg_r_1_26 ),
    .A1(tdc_inst_capt_out_26 ),
    .S(_0140_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_1 _0631_ (.A(_0133_),
    .B(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(_0148_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(tdc_inst_capt_reg_r_1_27 ),
    .A1(tdc_inst_capt_out_27 ),
    .S(_0140_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _0634_ (.A(_0133_),
    .B(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _0635_ (.A(_0150_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(tdc_inst_capt_reg_r_1_28 ),
    .A1(tdc_inst_capt_out_28 ),
    .S(_0140_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _0637_ (.A(_0133_),
    .B(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _0638_ (.A(_0152_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(tdc_inst_capt_reg_r_1_29 ),
    .A1(tdc_inst_capt_out_29 ),
    .S(_0140_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _0640_ (.A(_0133_),
    .B(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _0641_ (.A(_0154_),
    .X(_0032_));
 sky130_fd_sc_hd__clkbuf_2 _0642_ (.A(net2),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(tdc_inst_capt_reg_r_1_30 ),
    .A1(tdc_inst_capt_out_30 ),
    .S(_0140_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_1 _0644_ (.A(_0155_),
    .B(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _0645_ (.A(_0157_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(tdc_inst_capt_reg_r_1_31 ),
    .A1(tdc_inst_capt_out_31 ),
    .S(_0140_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_1 _0647_ (.A(_0155_),
    .B(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0159_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(tdc_inst_capt_reg_r_1_32 ),
    .A1(tdc_inst_capt_out_32 ),
    .S(_0140_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _0650_ (.A(_0155_),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(_0161_),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_4 _0652_ (.A(_0080_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0653_ (.A0(tdc_inst_capt_reg_r_1_33 ),
    .A1(tdc_inst_capt_out_33 ),
    .S(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _0654_ (.A(_0155_),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0655_ (.A(_0164_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0656_ (.A0(tdc_inst_capt_reg_r_1_34 ),
    .A1(tdc_inst_capt_out_34 ),
    .S(_0162_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_1 _0657_ (.A(_0155_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0658_ (.A(_0166_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(tdc_inst_capt_reg_r_1_35 ),
    .A1(tdc_inst_capt_out_35 ),
    .S(_0162_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _0660_ (.A(_0155_),
    .B(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0661_ (.A(_0168_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(tdc_inst_capt_reg_r_1_36 ),
    .A1(tdc_inst_capt_out_36 ),
    .S(_0162_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _0663_ (.A(_0155_),
    .B(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0170_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0665_ (.A0(tdc_inst_capt_reg_r_1_37 ),
    .A1(tdc_inst_capt_out_37 ),
    .S(_0162_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _0666_ (.A(_0155_),
    .B(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _0667_ (.A(_0172_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0668_ (.A0(tdc_inst_capt_reg_r_1_38 ),
    .A1(tdc_inst_capt_out_38 ),
    .S(_0162_),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _0669_ (.A(_0155_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_1 _0670_ (.A(_0174_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0671_ (.A0(tdc_inst_capt_reg_r_1_39 ),
    .A1(tdc_inst_capt_out_39 ),
    .S(_0162_),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _0672_ (.A(_0155_),
    .B(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_1 _0673_ (.A(_0176_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_2 _0674_ (.A(net2),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _0675_ (.A0(tdc_inst_capt_reg_r_1_40 ),
    .A1(tdc_inst_capt_out_40 ),
    .S(_0162_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _0676_ (.A(_0177_),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0677_ (.A(_0179_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(tdc_inst_capt_reg_r_1_41 ),
    .A1(tdc_inst_capt_out_41 ),
    .S(_0162_),
    .X(_0180_));
 sky130_fd_sc_hd__and2_1 _0679_ (.A(_0177_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(_0181_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0681_ (.A0(tdc_inst_capt_reg_r_1_42 ),
    .A1(tdc_inst_capt_out_42 ),
    .S(_0162_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_1 _0682_ (.A(_0177_),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _0683_ (.A(_0183_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _0684_ (.A(_0080_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _0685_ (.A0(tdc_inst_capt_reg_r_1_43 ),
    .A1(tdc_inst_capt_out_43 ),
    .S(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _0686_ (.A(_0177_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0687_ (.A(_0186_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(tdc_inst_capt_reg_r_1_44 ),
    .A1(tdc_inst_capt_out_44 ),
    .S(_0184_),
    .X(_0187_));
 sky130_fd_sc_hd__and2_1 _0689_ (.A(_0177_),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _0690_ (.A(_0188_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(tdc_inst_capt_reg_r_1_45 ),
    .A1(tdc_inst_capt_out_45 ),
    .S(_0184_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _0692_ (.A(_0177_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _0693_ (.A(_0190_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(tdc_inst_capt_reg_r_1_46 ),
    .A1(tdc_inst_capt_out_46 ),
    .S(_0184_),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _0695_ (.A(_0177_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0696_ (.A(_0192_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(tdc_inst_capt_reg_r_1_47 ),
    .A1(tdc_inst_capt_out_47 ),
    .S(_0184_),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _0698_ (.A(_0177_),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _0699_ (.A(_0194_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(tdc_inst_capt_reg_r_1_48 ),
    .A1(tdc_inst_capt_out_48 ),
    .S(_0184_),
    .X(_0195_));
 sky130_fd_sc_hd__and2_1 _0701_ (.A(_0177_),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _0702_ (.A(_0196_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(tdc_inst_capt_reg_r_1_49 ),
    .A1(tdc_inst_capt_out_49 ),
    .S(_0184_),
    .X(_0197_));
 sky130_fd_sc_hd__and2_1 _0704_ (.A(_0177_),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _0705_ (.A(_0198_),
    .X(_0052_));
 sky130_fd_sc_hd__buf_2 _0706_ (.A(net2),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(tdc_inst_capt_reg_r_1_50 ),
    .A1(tdc_inst_capt_out_50 ),
    .S(_0184_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(_0199_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0201_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(tdc_inst_capt_reg_r_1_51 ),
    .A1(tdc_inst_capt_out_51 ),
    .S(_0184_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(_0199_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0203_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(tdc_inst_capt_reg_r_1_52 ),
    .A1(tdc_inst_capt_out_52 ),
    .S(_0184_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _0714_ (.A(_0199_),
    .B(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _0715_ (.A(_0205_),
    .X(_0055_));
 sky130_fd_sc_hd__clkbuf_4 _0716_ (.A(_0080_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(tdc_inst_capt_reg_r_1_53 ),
    .A1(tdc_inst_capt_out_53 ),
    .S(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__and2_1 _0718_ (.A(_0199_),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _0719_ (.A(_0208_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(tdc_inst_capt_reg_r_1_54 ),
    .A1(tdc_inst_capt_out_54 ),
    .S(_0206_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _0721_ (.A(_0199_),
    .B(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _0722_ (.A(_0210_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(tdc_inst_capt_reg_r_1_55 ),
    .A1(tdc_inst_capt_out_55 ),
    .S(_0206_),
    .X(_0211_));
 sky130_fd_sc_hd__and2_1 _0724_ (.A(_0199_),
    .B(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _0725_ (.A(_0212_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(tdc_inst_capt_reg_r_1_56 ),
    .A1(tdc_inst_capt_out_56 ),
    .S(_0206_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(_0199_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _0728_ (.A(_0214_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(tdc_inst_capt_reg_r_1_57 ),
    .A1(tdc_inst_capt_out_57 ),
    .S(_0206_),
    .X(_0215_));
 sky130_fd_sc_hd__and2_1 _0730_ (.A(_0199_),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _0731_ (.A(_0216_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(tdc_inst_capt_reg_r_1_58 ),
    .A1(tdc_inst_capt_out_58 ),
    .S(_0206_),
    .X(_0217_));
 sky130_fd_sc_hd__and2_1 _0733_ (.A(_0199_),
    .B(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _0734_ (.A(_0218_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(tdc_inst_capt_reg_r_1_59 ),
    .A1(tdc_inst_capt_out_59 ),
    .S(_0206_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_1 _0736_ (.A(_0199_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0220_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(tdc_inst_capt_reg_r_1_60 ),
    .A1(tdc_inst_capt_out_60 ),
    .S(_0206_),
    .X(_0221_));
 sky130_fd_sc_hd__and2_1 _0739_ (.A(_0077_),
    .B(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _0740_ (.A(_0222_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(tdc_inst_capt_reg_r_1_61 ),
    .A1(tdc_inst_capt_out_61 ),
    .S(_0206_),
    .X(_0223_));
 sky130_fd_sc_hd__and2_1 _0742_ (.A(_0077_),
    .B(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0224_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(tdc_inst_capt_reg_r_1_62 ),
    .A1(tdc_inst_capt_out_62 ),
    .S(_0206_),
    .X(_0225_));
 sky130_fd_sc_hd__and2_1 _0745_ (.A(_0077_),
    .B(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _0746_ (.A(_0226_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0747_ (.A0(tdc_inst_capt_reg_r_1_63 ),
    .A1(tdc_inst_capt_out_63 ),
    .S(_0080_),
    .X(_0227_));
 sky130_fd_sc_hd__and2_1 _0748_ (.A(_0077_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _0749_ (.A(_0228_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(tdc_inst_pc_inst_val_in ),
    .A1(tdc_inst_val_out_capt ),
    .S(_0080_),
    .X(_0229_));
 sky130_fd_sc_hd__and2_1 _0751_ (.A(_0077_),
    .B(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_1 _0752_ (.A(_0230_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_2 _0753_ (.A(_0081_),
    .X(_0231_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(tdc_inst_capt_reg_r_1_60 ),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(tdc_inst_capt_reg_r_1_42 ),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(tdc_inst_capt_reg_r_1_58 ),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(tdc_inst_capt_reg_r_1_53 ),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(tdc_inst_capt_reg_r_1_49 ),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _0759_ (.A(tdc_inst_capt_reg_r_1_63 ),
    .B(tdc_inst_capt_reg_r_1_41 ),
    .Y(_0237_));
 sky130_fd_sc_hd__or2_1 _0760_ (.A(tdc_inst_capt_reg_r_1_63 ),
    .B(tdc_inst_capt_reg_r_1_41 ),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_2 _0761_ (.A(_0237_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__xor2_4 _0762_ (.A(tdc_inst_capt_reg_r_1_55 ),
    .B(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(tdc_inst_capt_reg_r_1_7 ),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2_1 _0764_ (.A(tdc_inst_capt_reg_r_1_14 ),
    .B(tdc_inst_capt_reg_r_1_10 ),
    .Y(_0242_));
 sky130_fd_sc_hd__or2_1 _0765_ (.A(tdc_inst_capt_reg_r_1_14 ),
    .B(tdc_inst_capt_reg_r_1_10 ),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _0766_ (.A(_0242_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__xor2_2 _0767_ (.A(tdc_inst_capt_reg_r_1_35 ),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xnor2_2 _0768_ (.A(_0241_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__xor2_2 _0769_ (.A(_0240_),
    .B(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__xor2_2 _0770_ (.A(tdc_inst_capt_reg_r_1_28 ),
    .B(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__xnor2_2 _0771_ (.A(tdc_inst_capt_reg_r_1_11 ),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(tdc_inst_capt_reg_r_1_38 ),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(tdc_inst_capt_reg_r_1_26 ),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(tdc_inst_capt_reg_r_1_24 ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(tdc_inst_capt_reg_r_1_3 ),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(tdc_inst_capt_reg_r_1_0 ),
    .Y(_0254_));
 sky130_fd_sc_hd__xor2_2 _0777_ (.A(tdc_inst_capt_reg_r_1_2 ),
    .B(tdc_inst_capt_reg_r_1_1 ),
    .X(_0255_));
 sky130_fd_sc_hd__xnor2_2 _0778_ (.A(tdc_inst_capt_reg_r_1_6 ),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__xnor2_2 _0779_ (.A(_0254_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__xnor2_2 _0780_ (.A(_0253_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__xnor2_1 _0781_ (.A(_0252_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__xnor2_1 _0782_ (.A(_0251_),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__xnor2_1 _0783_ (.A(_0250_),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__xor2_1 _0784_ (.A(_0249_),
    .B(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _0785_ (.A(tdc_inst_capt_reg_r_1_47 ),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__or2_1 _0786_ (.A(tdc_inst_capt_reg_r_1_47 ),
    .B(_0262_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_2 _0787_ (.A(_0263_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__xnor2_2 _0788_ (.A(_0236_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(tdc_inst_capt_reg_r_1_34 ),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(tdc_inst_capt_reg_r_1_32 ),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_2 _0791_ (.A(tdc_inst_capt_reg_r_1_13 ),
    .B(tdc_inst_capt_reg_r_1_9 ),
    .Y(_0269_));
 sky130_fd_sc_hd__or2_1 _0792_ (.A(tdc_inst_capt_reg_r_1_13 ),
    .B(tdc_inst_capt_reg_r_1_9 ),
    .X(_0270_));
 sky130_fd_sc_hd__a21o_1 _0793_ (.A1(_0269_),
    .A2(_0270_),
    .B1(tdc_inst_capt_reg_r_1_5 ),
    .X(_0271_));
 sky130_fd_sc_hd__nand3_2 _0794_ (.A(tdc_inst_capt_reg_r_1_5 ),
    .B(_0269_),
    .C(_0270_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _0795_ (.A(_0271_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(tdc_inst_capt_reg_r_1_4 ),
    .Y(_0274_));
 sky130_fd_sc_hd__xor2_2 _0797_ (.A(tdc_inst_capt_reg_r_1_21 ),
    .B(tdc_inst_capt_reg_r_1_19 ),
    .X(_0275_));
 sky130_fd_sc_hd__xnor2_2 _0798_ (.A(tdc_inst_capt_reg_r_1_17 ),
    .B(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__xnor2_1 _0799_ (.A(_0274_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_1 _0800_ (.A(_0273_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0273_),
    .B(_0277_),
    .Y(_0279_));
 sky130_fd_sc_hd__and2_1 _0802_ (.A(_0278_),
    .B(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(tdc_inst_capt_reg_r_1_22 ),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(tdc_inst_capt_reg_r_1_8 ),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(tdc_inst_capt_reg_r_1_12 ),
    .Y(_0283_));
 sky130_fd_sc_hd__xor2_1 _0806_ (.A(tdc_inst_capt_reg_r_1_27 ),
    .B(tdc_inst_capt_reg_r_1_25 ),
    .X(_0284_));
 sky130_fd_sc_hd__xnor2_1 _0807_ (.A(tdc_inst_capt_reg_r_1_23 ),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__xnor2_1 _0808_ (.A(_0283_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__xnor2_1 _0809_ (.A(_0282_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__xnor2_1 _0810_ (.A(_0281_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__xor2_1 _0811_ (.A(_0280_),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _0812_ (.A(_0268_),
    .B(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_1 _0813_ (.A(_0268_),
    .B(_0289_),
    .Y(_0291_));
 sky130_fd_sc_hd__nand2_1 _0814_ (.A(_0290_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__xnor2_2 _0815_ (.A(_0267_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(tdc_inst_capt_reg_r_1_20 ),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(tdc_inst_capt_reg_r_1_33 ),
    .B(tdc_inst_capt_reg_r_1_31 ),
    .Y(_0295_));
 sky130_fd_sc_hd__or2_1 _0818_ (.A(tdc_inst_capt_reg_r_1_33 ),
    .B(tdc_inst_capt_reg_r_1_31 ),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _0819_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__xor2_2 _0820_ (.A(tdc_inst_capt_reg_r_1_29 ),
    .B(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(tdc_inst_capt_reg_r_1_16 ),
    .Y(_0299_));
 sky130_fd_sc_hd__xor2_2 _0822_ (.A(tdc_inst_capt_reg_r_1_44 ),
    .B(tdc_inst_capt_reg_r_1_40 ),
    .X(_0300_));
 sky130_fd_sc_hd__xnor2_2 _0823_ (.A(tdc_inst_capt_reg_r_1_36 ),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_2 _0824_ (.A(_0299_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__xor2_2 _0825_ (.A(_0298_),
    .B(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__xnor2_2 _0826_ (.A(tdc_inst_capt_reg_r_1_18 ),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__xnor2_2 _0827_ (.A(_0294_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0828_ (.A(tdc_inst_capt_reg_r_1_37 ),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(tdc_inst_capt_reg_r_1_39 ),
    .Y(_0307_));
 sky130_fd_sc_hd__xor2_2 _0830_ (.A(tdc_inst_capt_reg_r_1_50 ),
    .B(tdc_inst_capt_reg_r_1_48 ),
    .X(_0308_));
 sky130_fd_sc_hd__xnor2_2 _0831_ (.A(tdc_inst_capt_reg_r_1_46 ),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__xnor2_2 _0832_ (.A(_0307_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__xnor2_2 _0833_ (.A(_0306_),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(tdc_inst_capt_reg_r_1_57 ),
    .B(tdc_inst_capt_reg_r_1_54 ),
    .Y(_0312_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(tdc_inst_capt_reg_r_1_57 ),
    .B(tdc_inst_capt_reg_r_1_54 ),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _0836_ (.A(_0312_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__xor2_2 _0837_ (.A(tdc_inst_capt_reg_r_1_52 ),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(tdc_inst_capt_reg_r_1_43 ),
    .Y(_0316_));
 sky130_fd_sc_hd__xor2_2 _0839_ (.A(tdc_inst_capt_reg_r_1_62 ),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0317_));
 sky130_fd_sc_hd__xnor2_2 _0840_ (.A(tdc_inst_capt_reg_r_1_59 ),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__xnor2_2 _0841_ (.A(_0316_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__xor2_2 _0842_ (.A(_0315_),
    .B(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__xnor2_2 _0843_ (.A(tdc_inst_capt_reg_r_1_15 ),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__xor2_2 _0844_ (.A(_0311_),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__xnor2_2 _0845_ (.A(tdc_inst_capt_reg_r_1_30 ),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__xor2_2 _0846_ (.A(_0305_),
    .B(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__xnor2_2 _0847_ (.A(tdc_inst_capt_reg_r_1_45 ),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__xor2_2 _0848_ (.A(_0293_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__xnor2_2 _0849_ (.A(tdc_inst_capt_reg_r_1_51 ),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__xor2_2 _0850_ (.A(_0266_),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__xnor2_2 _0851_ (.A(tdc_inst_capt_reg_r_1_56 ),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__xnor2_2 _0852_ (.A(_0235_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xnor2_2 _0853_ (.A(_0234_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__xnor2_2 _0854_ (.A(_0233_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(_0232_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(_0232_),
    .B(_0332_),
    .X(_0334_));
 sky130_fd_sc_hd__o21ai_1 _0857_ (.A1(_0333_),
    .A2(_0334_),
    .B1(_0231_),
    .Y(_0335_));
 sky130_fd_sc_hd__o211a_1 _0858_ (.A1(_0231_),
    .A2(net35),
    .B1(_0078_),
    .C1(_0335_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _0859_ (.A(tdc_inst_capt_reg_r_1_28 ),
    .B(_0247_),
    .X(_0336_));
 sky130_fd_sc_hd__a21o_1 _0860_ (.A1(tdc_inst_capt_reg_r_1_11 ),
    .A2(_0248_),
    .B1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__o21ai_2 _0861_ (.A1(_0236_),
    .A2(_0265_),
    .B1(_0263_),
    .Y(_0338_));
 sky130_fd_sc_hd__or2_1 _0862_ (.A(_0250_),
    .B(_0260_),
    .X(_0339_));
 sky130_fd_sc_hd__o21a_1 _0863_ (.A1(_0249_),
    .A2(_0261_),
    .B1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_2 _0864_ (.A1(_0267_),
    .A2(_0292_),
    .B1(_0290_),
    .Y(_0341_));
 sky130_fd_sc_hd__a21bo_1 _0865_ (.A1(tdc_inst_capt_reg_r_1_55 ),
    .A2(_0238_),
    .B1_N(_0237_),
    .X(_0342_));
 sky130_fd_sc_hd__a21bo_1 _0866_ (.A1(tdc_inst_capt_reg_r_1_35 ),
    .A2(_0243_),
    .B1_N(_0242_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _0867_ (.A(_0241_),
    .B(_0245_),
    .X(_0344_));
 sky130_fd_sc_hd__o21a_1 _0868_ (.A1(_0240_),
    .A2(_0246_),
    .B1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__xnor2_2 _0869_ (.A(_0343_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__xor2_2 _0870_ (.A(_0342_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _0871_ (.A(_0254_),
    .B(_0256_),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_2 _0872_ (.A1(_0253_),
    .A2(_0257_),
    .B1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__o21ai_1 _0873_ (.A1(_0274_),
    .A2(_0276_),
    .B1(_0278_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _0874_ (.A(tdc_inst_capt_reg_r_1_2 ),
    .B(tdc_inst_capt_reg_r_1_1 ),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _0875_ (.A(tdc_inst_capt_reg_r_1_6 ),
    .B(_0255_),
    .Y(_0352_));
 sky130_fd_sc_hd__a22oi_4 _0876_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0269_),
    .B2(_0272_),
    .Y(_0353_));
 sky130_fd_sc_hd__and4_1 _0877_ (.A(_0351_),
    .B(_0352_),
    .C(_0269_),
    .D(_0272_),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_1 _0878_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__xnor2_1 _0879_ (.A(_0350_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__xor2_2 _0880_ (.A(_0349_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _0881_ (.A(_0252_),
    .B(_0258_),
    .X(_0358_));
 sky130_fd_sc_hd__o21a_1 _0882_ (.A1(_0251_),
    .A2(_0259_),
    .B1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__xor2_2 _0883_ (.A(_0357_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__xnor2_2 _0884_ (.A(_0347_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__xnor2_2 _0885_ (.A(_0341_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__xnor2_2 _0886_ (.A(_0340_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(_0281_),
    .B(_0287_),
    .X(_0364_));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(_0288_),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _0889_ (.A(_0280_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _0890_ (.A(tdc_inst_capt_reg_r_1_18 ),
    .B(_0303_),
    .Y(_0367_));
 sky130_fd_sc_hd__o21a_1 _0891_ (.A1(_0294_),
    .A2(_0304_),
    .B1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _0892_ (.A(tdc_inst_capt_reg_r_1_21 ),
    .B(tdc_inst_capt_reg_r_1_19 ),
    .X(_0369_));
 sky130_fd_sc_hd__a21oi_1 _0893_ (.A1(tdc_inst_capt_reg_r_1_17 ),
    .A2(_0275_),
    .B1(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21boi_1 _0894_ (.A1(tdc_inst_capt_reg_r_1_29 ),
    .A2(_0296_),
    .B1_N(_0295_),
    .Y(_0371_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(tdc_inst_capt_reg_r_1_27 ),
    .B(tdc_inst_capt_reg_r_1_25 ),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _0896_ (.A1(tdc_inst_capt_reg_r_1_23 ),
    .A2(_0284_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__or2_1 _0897_ (.A(_0371_),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _0898_ (.A(_0371_),
    .B(_0373_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _0899_ (.A(_0374_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__or2_1 _0900_ (.A(_0283_),
    .B(_0285_),
    .X(_0377_));
 sky130_fd_sc_hd__o21a_1 _0901_ (.A1(_0282_),
    .A2(_0286_),
    .B1(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__xnor2_1 _0902_ (.A(_0376_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__xnor2_1 _0903_ (.A(_0370_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__xnor2_1 _0904_ (.A(_0368_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__a21o_1 _0905_ (.A1(_0364_),
    .A2(_0366_),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nand3_1 _0906_ (.A(_0364_),
    .B(_0366_),
    .C(_0381_),
    .Y(_0383_));
 sky130_fd_sc_hd__and2_2 _0907_ (.A(_0382_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__or2_1 _0908_ (.A(_0299_),
    .B(_0301_),
    .X(_0385_));
 sky130_fd_sc_hd__o21a_1 _0909_ (.A1(_0298_),
    .A2(_0302_),
    .B1(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _0910_ (.A(_0307_),
    .B(_0309_),
    .X(_0387_));
 sky130_fd_sc_hd__o21a_1 _0911_ (.A1(_0306_),
    .A2(_0310_),
    .B1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _0912_ (.A(tdc_inst_capt_reg_r_1_44 ),
    .B(tdc_inst_capt_reg_r_1_40 ),
    .X(_0389_));
 sky130_fd_sc_hd__a21oi_2 _0913_ (.A1(tdc_inst_capt_reg_r_1_36 ),
    .A2(_0300_),
    .B1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__xor2_2 _0914_ (.A(_0388_),
    .B(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__xnor2_2 _0915_ (.A(_0386_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21bo_2 _0916_ (.A1(tdc_inst_capt_reg_r_1_52 ),
    .A2(_0313_),
    .B1_N(_0312_),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(tdc_inst_capt_reg_r_1_50 ),
    .B(tdc_inst_capt_reg_r_1_48 ),
    .X(_0394_));
 sky130_fd_sc_hd__a21o_1 _0918_ (.A1(tdc_inst_capt_reg_r_1_46 ),
    .A2(_0308_),
    .B1(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__xor2_4 _0919_ (.A(_0393_),
    .B(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _0920_ (.A(tdc_inst_capt_reg_r_1_62 ),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0397_));
 sky130_fd_sc_hd__a21o_2 _0921_ (.A1(tdc_inst_capt_reg_r_1_59 ),
    .A2(_0317_),
    .B1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _0922_ (.A(_0316_),
    .B(_0318_),
    .X(_0399_));
 sky130_fd_sc_hd__o21a_2 _0923_ (.A1(_0315_),
    .A2(_0319_),
    .B1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__xnor2_4 _0924_ (.A(_0398_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_2 _0925_ (.A(_0396_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _0926_ (.A(tdc_inst_capt_reg_r_1_15 ),
    .B(_0320_),
    .Y(_0403_));
 sky130_fd_sc_hd__o21a_1 _0927_ (.A1(_0311_),
    .A2(_0321_),
    .B1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__xor2_2 _0928_ (.A(_0402_),
    .B(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__xnor2_2 _0929_ (.A(_0392_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _0930_ (.A(tdc_inst_capt_reg_r_1_30 ),
    .B(_0322_),
    .Y(_0407_));
 sky130_fd_sc_hd__o21ai_2 _0931_ (.A1(_0305_),
    .A2(_0323_),
    .B1(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__xnor2_2 _0932_ (.A(_0406_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_2 _0933_ (.A(_0384_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _0934_ (.A(tdc_inst_capt_reg_r_1_45 ),
    .B(_0324_),
    .Y(_0411_));
 sky130_fd_sc_hd__o21ai_2 _0935_ (.A1(_0293_),
    .A2(_0325_),
    .B1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__xnor2_2 _0936_ (.A(_0410_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__xnor2_2 _0937_ (.A(_0363_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(tdc_inst_capt_reg_r_1_51 ),
    .B(_0326_),
    .Y(_0415_));
 sky130_fd_sc_hd__o21a_1 _0939_ (.A1(_0266_),
    .A2(_0327_),
    .B1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__xor2_2 _0940_ (.A(_0414_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__xnor2_2 _0941_ (.A(_0338_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _0942_ (.A(tdc_inst_capt_reg_r_1_56 ),
    .B(_0328_),
    .Y(_0419_));
 sky130_fd_sc_hd__o21a_1 _0943_ (.A1(_0235_),
    .A2(_0329_),
    .B1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__xnor2_1 _0944_ (.A(_0418_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__xor2_1 _0945_ (.A(_0337_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_1 _0946_ (.A(_0234_),
    .B(_0330_),
    .X(_0423_));
 sky130_fd_sc_hd__o21a_1 _0947_ (.A1(_0233_),
    .A2(_0331_),
    .B1(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__xor2_1 _0948_ (.A(_0422_),
    .B(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__xnor2_1 _0949_ (.A(_0333_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__nand2_1 _0950_ (.A(_0231_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__o211a_1 _0951_ (.A1(_0231_),
    .A2(uo_out[1]),
    .B1(_0078_),
    .C1(_0427_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _0952_ (.A(_0418_),
    .B(_0420_),
    .X(_0428_));
 sky130_fd_sc_hd__or2b_1 _0953_ (.A(_0421_),
    .B_N(_0337_),
    .X(_0429_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(_0345_),
    .Y(_0430_));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(_0342_),
    .B(_0346_),
    .X(_0431_));
 sky130_fd_sc_hd__a21o_1 _0956_ (.A1(_0343_),
    .A2(_0430_),
    .B1(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__or2b_1 _0957_ (.A(_0361_),
    .B_N(_0341_),
    .X(_0433_));
 sky130_fd_sc_hd__or2b_1 _0958_ (.A(_0340_),
    .B_N(_0362_),
    .X(_0434_));
 sky130_fd_sc_hd__nand2_1 _0959_ (.A(_0433_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _0960_ (.A(_0357_),
    .B(_0359_),
    .Y(_0436_));
 sky130_fd_sc_hd__a21o_1 _0961_ (.A1(_0347_),
    .A2(_0360_),
    .B1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__o21ai_1 _0962_ (.A1(_0368_),
    .A2(_0380_),
    .B1(_0382_),
    .Y(_0438_));
 sky130_fd_sc_hd__and2b_1 _0963_ (.A_N(_0356_),
    .B(_0349_),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _0964_ (.A1(_0350_),
    .A2(_0355_),
    .B1(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__xnor2_2 _0965_ (.A(_0353_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__xor2_1 _0966_ (.A(_0438_),
    .B(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__xor2_1 _0967_ (.A(_0437_),
    .B(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__or2_1 _0968_ (.A(_0376_),
    .B(_0378_),
    .X(_0444_));
 sky130_fd_sc_hd__o21ai_1 _0969_ (.A1(_0370_),
    .A2(_0379_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__and2b_1 _0970_ (.A_N(_0386_),
    .B(_0391_),
    .X(_0446_));
 sky130_fd_sc_hd__o21ba_1 _0971_ (.A1(_0388_),
    .A2(_0390_),
    .B1_N(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__xnor2_1 _0972_ (.A(_0374_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__xnor2_1 _0973_ (.A(_0445_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__nor2_1 _0974_ (.A(_0402_),
    .B(_0404_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21oi_1 _0975_ (.A1(_0392_),
    .A2(_0405_),
    .B1(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__and2_1 _0976_ (.A(_0393_),
    .B(_0395_),
    .X(_0452_));
 sky130_fd_sc_hd__inv_2 _0977_ (.A(_0398_),
    .Y(_0453_));
 sky130_fd_sc_hd__nor2_1 _0978_ (.A(_0453_),
    .B(_0400_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand2_2 _0979_ (.A(_0452_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__or2_1 _0980_ (.A(_0452_),
    .B(_0454_),
    .X(_0456_));
 sky130_fd_sc_hd__a22oi_4 _0981_ (.A1(_0396_),
    .A2(_0401_),
    .B1(_0455_),
    .B2(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__xor2_1 _0982_ (.A(_0451_),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__xnor2_1 _0983_ (.A(_0449_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__or2b_1 _0984_ (.A(_0406_),
    .B_N(_0408_),
    .X(_0460_));
 sky130_fd_sc_hd__a21boi_2 _0985_ (.A1(_0384_),
    .A2(_0409_),
    .B1_N(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__xor2_1 _0986_ (.A(_0459_),
    .B(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__xnor2_1 _0987_ (.A(_0443_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__and2b_1 _0988_ (.A_N(_0410_),
    .B(_0412_),
    .X(_0464_));
 sky130_fd_sc_hd__a21oi_1 _0989_ (.A1(_0363_),
    .A2(_0413_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__xnor2_1 _0990_ (.A(_0463_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__xor2_1 _0991_ (.A(_0435_),
    .B(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__nor2_1 _0992_ (.A(_0414_),
    .B(_0416_),
    .Y(_0468_));
 sky130_fd_sc_hd__a21oi_1 _0993_ (.A1(_0338_),
    .A2(_0417_),
    .B1(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__xor2_1 _0994_ (.A(_0467_),
    .B(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__xnor2_1 _0995_ (.A(_0432_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__a21o_1 _0996_ (.A1(_0428_),
    .A2(_0429_),
    .B1(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__nand3_1 _0997_ (.A(_0428_),
    .B(_0429_),
    .C(_0471_),
    .Y(_0473_));
 sky130_fd_sc_hd__and2_1 _0998_ (.A(_0472_),
    .B(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _0999_ (.A(_0422_),
    .B(_0424_),
    .Y(_0475_));
 sky130_fd_sc_hd__a21o_1 _1000_ (.A1(_0333_),
    .A2(_0425_),
    .B1(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0474_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__or2_1 _1002_ (.A(_0474_),
    .B(_0476_),
    .X(_0478_));
 sky130_fd_sc_hd__a21bo_1 _1003_ (.A1(_0477_),
    .A2(_0478_),
    .B1_N(_0231_),
    .X(_0479_));
 sky130_fd_sc_hd__o211a_1 _1004_ (.A1(_0231_),
    .A2(net37),
    .B1(_0078_),
    .C1(_0479_),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _1005_ (.A(_0467_),
    .B(_0469_),
    .X(_0480_));
 sky130_fd_sc_hd__nand2_1 _1006_ (.A(_0432_),
    .B(_0470_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0438_),
    .B(_0441_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21bo_1 _1008_ (.A1(_0437_),
    .A2(_0442_),
    .B1_N(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__nand2_1 _1009_ (.A(_0353_),
    .B(_0439_),
    .Y(_0484_));
 sky130_fd_sc_hd__or2b_1 _1010_ (.A(_0448_),
    .B_N(_0445_),
    .X(_0485_));
 sky130_fd_sc_hd__o21a_1 _1011_ (.A1(_0374_),
    .A2(_0447_),
    .B1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(_0484_),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__nand2_1 _1013_ (.A(_0484_),
    .B(_0486_),
    .Y(_0488_));
 sky130_fd_sc_hd__and2_1 _1014_ (.A(_0487_),
    .B(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nor2_1 _1015_ (.A(_0451_),
    .B(_0457_),
    .Y(_0490_));
 sky130_fd_sc_hd__a21oi_1 _1016_ (.A1(_0449_),
    .A2(_0458_),
    .B1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _1017_ (.A(_0455_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _1018_ (.A(_0455_),
    .B(_0491_),
    .Y(_0493_));
 sky130_fd_sc_hd__and2_1 _1019_ (.A(_0492_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__xnor2_1 _1020_ (.A(_0489_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__nor2_1 _1021_ (.A(_0459_),
    .B(_0461_),
    .Y(_0496_));
 sky130_fd_sc_hd__a21oi_1 _1022_ (.A1(_0443_),
    .A2(_0462_),
    .B1(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__xnor2_1 _1023_ (.A(_0495_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__xor2_1 _1024_ (.A(_0483_),
    .B(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__or2b_1 _1025_ (.A(_0466_),
    .B_N(_0435_),
    .X(_0500_));
 sky130_fd_sc_hd__o21a_1 _1026_ (.A1(_0463_),
    .A2(_0465_),
    .B1(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__xnor2_1 _1027_ (.A(_0499_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__and3_1 _1028_ (.A(_0480_),
    .B(_0481_),
    .C(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__a21o_1 _1029_ (.A1(_0480_),
    .A2(_0481_),
    .B1(_0502_),
    .X(_0504_));
 sky130_fd_sc_hd__and2b_1 _1030_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__a21o_1 _1031_ (.A1(_0472_),
    .A2(_0477_),
    .B1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _1032_ (.A(_0081_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__a31o_1 _1033_ (.A1(_0472_),
    .A2(_0477_),
    .A3(_0505_),
    .B1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__o211a_1 _1034_ (.A1(_0231_),
    .A2(net38),
    .B1(_0078_),
    .C1(_0508_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _1035_ (.A(_0499_),
    .B(_0501_),
    .X(_0509_));
 sky130_fd_sc_hd__and2b_1 _1036_ (.A_N(_0498_),
    .B(_0483_),
    .X(_0510_));
 sky130_fd_sc_hd__o21bai_1 _1037_ (.A1(_0495_),
    .A2(_0497_),
    .B1_N(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21bo_1 _1038_ (.A1(_0489_),
    .A2(_0494_),
    .B1_N(_0492_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(_0492_),
    .A1(_0512_),
    .S(_0487_),
    .X(_0513_));
 sky130_fd_sc_hd__xnor2_1 _1040_ (.A(_0511_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _1041_ (.A(_0509_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__and2_1 _1042_ (.A(_0509_),
    .B(_0514_),
    .X(_0516_));
 sky130_fd_sc_hd__nor2_1 _1043_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__a21oi_1 _1044_ (.A1(_0472_),
    .A2(_0504_),
    .B1(_0503_),
    .Y(_0518_));
 sky130_fd_sc_hd__a31o_1 _1045_ (.A1(_0474_),
    .A2(_0476_),
    .A3(_0505_),
    .B1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__xnor2_1 _1046_ (.A(_0517_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _1047_ (.A(_0231_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__o211a_1 _1048_ (.A1(_0231_),
    .A2(net34),
    .B1(_0078_),
    .C1(_0521_),
    .X(_0072_));
 sky130_fd_sc_hd__and2b_1 _1049_ (.A_N(_0081_),
    .B(uo_out[5]),
    .X(_0522_));
 sky130_fd_sc_hd__o2bb2a_1 _1050_ (.A1_N(_0511_),
    .A2_N(_0513_),
    .B1(_0487_),
    .B2(_0492_),
    .X(_0523_));
 sky130_fd_sc_hd__a21oi_1 _1051_ (.A1(_0517_),
    .A2(_0519_),
    .B1(_0515_),
    .Y(_0524_));
 sky130_fd_sc_hd__o21ai_1 _1052_ (.A1(_0523_),
    .A2(_0524_),
    .B1(_0081_),
    .Y(_0525_));
 sky130_fd_sc_hd__a21oi_1 _1053_ (.A1(_0523_),
    .A2(_0524_),
    .B1(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__o21a_1 _1054_ (.A1(_0522_),
    .A2(_0526_),
    .B1(_0078_),
    .X(_0073_));
 sky130_fd_sc_hd__o211a_1 _1055_ (.A1(_0231_),
    .A2(net36),
    .B1(_0078_),
    .C1(_0525_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(tdc_inst_pc_inst_val_out ),
    .A1(tdc_inst_pc_inst_val_in ),
    .S(_0080_),
    .X(_0527_));
 sky130_fd_sc_hd__and2_1 _1057_ (.A(_0077_),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _1058_ (.A(_0528_),
    .X(_0075_));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_1_0__leaf_ui_in[0]),
    .D(_0000_),
    .Q(tdc_inst_pg_pg_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_1_1__leaf_ui_in[0]),
    .D(_0001_),
    .Q(tdc_inst_pg_val_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0002_),
    .Q(tdc_inst_val_out_capt ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0003_),
    .Q(tdc_inst_capt_reg_r_1_0 ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(_0004_),
    .Q(tdc_inst_capt_reg_r_1_1 ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0005_),
    .Q(tdc_inst_capt_reg_r_1_2 ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0006_),
    .Q(tdc_inst_capt_reg_r_1_3 ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0007_),
    .Q(tdc_inst_capt_reg_r_1_4 ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(_0008_),
    .Q(tdc_inst_capt_reg_r_1_5 ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0009_),
    .Q(tdc_inst_capt_reg_r_1_6 ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0010_),
    .Q(tdc_inst_capt_reg_r_1_7 ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0011_),
    .Q(tdc_inst_capt_reg_r_1_8 ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(_0012_),
    .Q(tdc_inst_capt_reg_r_1_9 ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0013_),
    .Q(tdc_inst_capt_reg_r_1_10 ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0014_),
    .Q(tdc_inst_capt_reg_r_1_11 ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0015_),
    .Q(tdc_inst_capt_reg_r_1_12 ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0016_),
    .Q(tdc_inst_capt_reg_r_1_13 ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0017_),
    .Q(tdc_inst_capt_reg_r_1_14 ));
 sky130_fd_sc_hd__dfxtp_2 _1077_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0018_),
    .Q(tdc_inst_capt_reg_r_1_15 ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0019_),
    .Q(tdc_inst_capt_reg_r_1_16 ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0020_),
    .Q(tdc_inst_capt_reg_r_1_17 ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0021_),
    .Q(tdc_inst_capt_reg_r_1_18 ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0022_),
    .Q(tdc_inst_capt_reg_r_1_19 ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0023_),
    .Q(tdc_inst_capt_reg_r_1_20 ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0024_),
    .Q(tdc_inst_capt_reg_r_1_21 ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0025_),
    .Q(tdc_inst_capt_reg_r_1_22 ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0026_),
    .Q(tdc_inst_capt_reg_r_1_23 ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0027_),
    .Q(tdc_inst_capt_reg_r_1_24 ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0028_),
    .Q(tdc_inst_capt_reg_r_1_25 ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0029_),
    .Q(tdc_inst_capt_reg_r_1_26 ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(_0030_),
    .Q(tdc_inst_capt_reg_r_1_27 ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0031_),
    .Q(tdc_inst_capt_reg_r_1_28 ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0032_),
    .Q(tdc_inst_capt_reg_r_1_29 ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0033_),
    .Q(tdc_inst_capt_reg_r_1_30 ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0034_),
    .Q(tdc_inst_capt_reg_r_1_31 ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0035_),
    .Q(tdc_inst_capt_reg_r_1_32 ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0036_),
    .Q(tdc_inst_capt_reg_r_1_33 ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0037_),
    .Q(tdc_inst_capt_reg_r_1_34 ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0038_),
    .Q(tdc_inst_capt_reg_r_1_35 ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0039_),
    .Q(tdc_inst_capt_reg_r_1_36 ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0040_),
    .Q(tdc_inst_capt_reg_r_1_37 ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0041_),
    .Q(tdc_inst_capt_reg_r_1_38 ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0042_),
    .Q(tdc_inst_capt_reg_r_1_39 ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0043_),
    .Q(tdc_inst_capt_reg_r_1_40 ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0044_),
    .Q(tdc_inst_capt_reg_r_1_41 ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0045_),
    .Q(tdc_inst_capt_reg_r_1_42 ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0046_),
    .Q(tdc_inst_capt_reg_r_1_43 ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0047_),
    .Q(tdc_inst_capt_reg_r_1_44 ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0048_),
    .Q(tdc_inst_capt_reg_r_1_45 ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0049_),
    .Q(tdc_inst_capt_reg_r_1_46 ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0050_),
    .Q(tdc_inst_capt_reg_r_1_47 ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0051_),
    .Q(tdc_inst_capt_reg_r_1_48 ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0052_),
    .Q(tdc_inst_capt_reg_r_1_49 ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0053_),
    .Q(tdc_inst_capt_reg_r_1_50 ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0054_),
    .Q(tdc_inst_capt_reg_r_1_51 ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0055_),
    .Q(tdc_inst_capt_reg_r_1_52 ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0056_),
    .Q(tdc_inst_capt_reg_r_1_53 ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0057_),
    .Q(tdc_inst_capt_reg_r_1_54 ));
 sky130_fd_sc_hd__dfxtp_2 _1117_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0058_),
    .Q(tdc_inst_capt_reg_r_1_55 ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0059_),
    .Q(tdc_inst_capt_reg_r_1_56 ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0060_),
    .Q(tdc_inst_capt_reg_r_1_57 ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0061_),
    .Q(tdc_inst_capt_reg_r_1_58 ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0062_),
    .Q(tdc_inst_capt_reg_r_1_59 ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0063_),
    .Q(tdc_inst_capt_reg_r_1_60 ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0064_),
    .Q(tdc_inst_capt_reg_r_1_61 ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(_0065_),
    .Q(tdc_inst_capt_reg_r_1_62 ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0066_),
    .Q(tdc_inst_capt_reg_r_1_63 ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0067_),
    .Q(tdc_inst_pc_inst_val_in ));
 sky130_fd_sc_hd__dfxtp_4 _1127_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0068_),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_4 _1128_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0069_),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_4 _1129_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0070_),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_4 _1130_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0071_),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_4 _1131_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0072_),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_4 _1132_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0073_),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_4 _1133_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0074_),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0075_),
    .Q(tdc_inst_pc_inst_val_out ));
 sky130_fd_sc_hd__buf_2 _1151_ (.A(tdc_inst_dl_inst_dl_genblk_dl_c_64 ),
    .X(tdc_inst_dl_inst_dl_genblk_dl_co ));
 sky130_fd_sc_hd__buf_2 _1152_ (.A(tdc_inst_dl_inst_dl_genblk_dl_c_0 ),
    .X(tdc_inst_pg_out ));
 sky130_fd_sc_hd__clkbuf_4 _1153_ (.A(tdc_inst_pc_inst_val_out ),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_ui_in_0  (.A(ui_in[0]),
    .X(clknet_0_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_ui_in_1  (.A(ui_in[1]),
    .X(clknet_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_ui_in_0  (.A(clknet_0_ui_in[0]),
    .X(clknet_1_0__leaf_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_ui_in_0  (.A(clknet_0_ui_in[0]),
    .X(clknet_1_1__leaf_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_0_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_10_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_11_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_12_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_13_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_14_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_15_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_1_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_2_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_3_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_4_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_5_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_6_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_7_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_8_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_9_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net16),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(net16),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net16),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net16),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net16),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(net16),
    .X(net8));
 sky130_fd_sc_hd__buf_2 fanout9 (.A(net16),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(tdc_inst_pg_val_r_out ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(uo_out[4]),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(uo_out[0]),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(uo_out[6]),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(uo_out[2]),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(uo_out[3]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input1 (.A(ena),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_0_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_0 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_0 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_10_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_10 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_10 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_11_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_11 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_11 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_12_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_12 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_12 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_13_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_13 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_13 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_14_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_14 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_14 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_15_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_15 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_15 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_16_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_16 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_16 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_17_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_17 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_17 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_18_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_18 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_18 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_19_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_19 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_19 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_1_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_1 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_1 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_20_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_20 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_20 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_21_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_21 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_21 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_22_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_22 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_22 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_23_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_23 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_23 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_24_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_24 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_24 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_25_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_25 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_25 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_26_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_26 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_26 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_27_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_27 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_27 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_28_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_28 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_28 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_29_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_29 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_29 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_2_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_2 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_2 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_30_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_30 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_30 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_31_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_31 ),
    .DE(net12),
    .Q(tdc_inst_capt_out_31 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_32_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_32 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_32 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_33_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_33 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_33 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_34_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_34 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_34 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_35_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_35 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_35 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_36_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_36 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_36 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_37_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_37 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_37 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_38_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_38 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_38 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_39_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_39 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_39 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_3_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_3 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_3 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_40_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_40 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_40 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_41_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_41 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_41 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_42_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_42 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_42 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_43_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_43 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_43 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_44_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_44 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_44 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_45_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_45 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_45 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_46_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_46 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_46 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_47_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_47 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_47 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_48_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_48 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_48 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_49_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_49 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_49 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_4_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_4 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_4 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_50_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_50 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_50 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_51_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_51 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_51 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_52_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_52 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_52 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_53_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_53 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_53 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_54_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_54 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_54 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_55_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_55 ),
    .DE(net9),
    .Q(tdc_inst_capt_out_55 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_56_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_56 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_56 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_57_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_57 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_57 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_58_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_58 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_58 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_59_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_59 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_59 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_5_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_5 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_5 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_60_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_60 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_60 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_61_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_61 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_61 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_62_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_62 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_62 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_63_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_63 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_63 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_6_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_6 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_6 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_7_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_7 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_7 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_8_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_8 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_8 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_9_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_capt_D_9 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_9 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_0_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_0 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_10_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_10 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_11_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_11 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_12_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_12 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_13_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_13 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_14_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_14 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_15_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_15 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_16_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_16 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_17_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_17 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_18_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_18 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_19_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_19 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_1_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_1 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_20_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_20 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_21_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_21 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_22_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_22 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_23_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_23 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_24_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_24 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_25_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_25 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_26_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_26 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_27_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_27 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_28_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_28 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_29_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_29 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_2_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_2 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_30_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_30 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_31_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_31 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_32_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_32 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_33_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_33 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_34_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_34 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_35_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_35 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_36_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_36 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_37_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_37 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_38_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_38 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_39_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_39 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_3_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_3 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_40_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_40 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_41_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_41 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_42_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_42 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_43_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_43 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_44_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_44 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_45_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_45 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_46_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_46 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_47_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_47 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_48_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_48 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_49_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_49 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_4_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_4 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_50_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_50 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_51_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_51 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_52_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_52 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_53_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_53 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_54_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_54 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_55_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_55 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_56_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_56 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_57_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_57 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_58_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_58 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_59_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_59 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_5_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_5 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_60_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_60 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_61_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_61 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_62_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_62 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_63_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_63 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_6_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_6 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_7_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_7 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_8_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_8 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_9_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_9 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_0_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_0 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_0 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_0 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_1 ),
    .SUM(tdc_inst_dl_capt_D_0 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_10_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_10 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_10 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_10 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_11 ),
    .SUM(tdc_inst_dl_capt_D_10 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_11_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_11 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_11 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_11 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_12 ),
    .SUM(tdc_inst_dl_capt_D_11 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_12_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_12 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_12 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_12 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_13 ),
    .SUM(tdc_inst_dl_capt_D_12 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_13_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_13 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_13 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_13 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_14 ),
    .SUM(tdc_inst_dl_capt_D_13 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_14_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_14 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_14 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_14 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_15 ),
    .SUM(tdc_inst_dl_capt_D_14 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_15_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_15 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_15 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_15 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_16 ),
    .SUM(tdc_inst_dl_capt_D_15 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_16_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_16 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_16 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_16 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_17 ),
    .SUM(tdc_inst_dl_capt_D_16 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_17_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_17 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_17 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_17 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_18 ),
    .SUM(tdc_inst_dl_capt_D_17 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_18_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_18 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_18 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_18 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_19 ),
    .SUM(tdc_inst_dl_capt_D_18 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_19_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_19 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_19 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_19 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_20 ),
    .SUM(tdc_inst_dl_capt_D_19 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_1_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_1 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_1 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_1 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_2 ),
    .SUM(tdc_inst_dl_capt_D_1 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_20_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_20 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_20 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_20 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_21 ),
    .SUM(tdc_inst_dl_capt_D_20 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_21_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_21 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_21 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_21 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_22 ),
    .SUM(tdc_inst_dl_capt_D_21 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_22_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_22 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_22 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_22 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_23 ),
    .SUM(tdc_inst_dl_capt_D_22 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_23_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_23 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_23 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_23 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_24 ),
    .SUM(tdc_inst_dl_capt_D_23 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_24_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_24 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_24 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_24 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_25 ),
    .SUM(tdc_inst_dl_capt_D_24 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_25_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_25 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_25 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_25 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_26 ),
    .SUM(tdc_inst_dl_capt_D_25 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_26_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_26 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_26 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_26 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_27 ),
    .SUM(tdc_inst_dl_capt_D_26 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_27_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_27 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_27 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_27 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_28 ),
    .SUM(tdc_inst_dl_capt_D_27 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_28_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_28 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_28 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_28 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_29 ),
    .SUM(tdc_inst_dl_capt_D_28 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_29_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_29 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_29 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_29 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_30 ),
    .SUM(tdc_inst_dl_capt_D_29 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_2_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_2 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_2 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_2 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_3 ),
    .SUM(tdc_inst_dl_capt_D_2 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_30_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_30 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_30 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_30 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_31 ),
    .SUM(tdc_inst_dl_capt_D_30 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_31_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_31 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_31 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_31 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_32 ),
    .SUM(tdc_inst_dl_capt_D_31 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_32_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_32 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_32 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_32 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_33 ),
    .SUM(tdc_inst_dl_capt_D_32 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_33_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_33 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_33 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_33 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_34 ),
    .SUM(tdc_inst_dl_capt_D_33 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_34_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_34 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_34 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_34 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_35 ),
    .SUM(tdc_inst_dl_capt_D_34 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_35_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_35 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_35 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_35 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_36 ),
    .SUM(tdc_inst_dl_capt_D_35 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_36_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_36 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_36 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_36 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_37 ),
    .SUM(tdc_inst_dl_capt_D_36 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_37_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_37 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_37 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_37 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_38 ),
    .SUM(tdc_inst_dl_capt_D_37 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_38_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_38 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_38 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_38 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_39 ),
    .SUM(tdc_inst_dl_capt_D_38 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_39_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_39 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_39 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_39 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_40 ),
    .SUM(tdc_inst_dl_capt_D_39 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_3_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_3 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_3 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_3 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_4 ),
    .SUM(tdc_inst_dl_capt_D_3 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_40_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_40 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_40 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_40 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_41 ),
    .SUM(tdc_inst_dl_capt_D_40 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_41_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_41 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_41 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_41 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_42 ),
    .SUM(tdc_inst_dl_capt_D_41 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_42_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_42 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_42 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_42 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_43 ),
    .SUM(tdc_inst_dl_capt_D_42 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_43_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_43 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_43 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_43 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_44 ),
    .SUM(tdc_inst_dl_capt_D_43 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_44_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_44 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_44 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_44 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_45 ),
    .SUM(tdc_inst_dl_capt_D_44 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_45_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_45 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_45 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_45 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_46 ),
    .SUM(tdc_inst_dl_capt_D_45 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_46_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_46 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_46 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_46 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_47 ),
    .SUM(tdc_inst_dl_capt_D_46 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_47_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_47 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_47 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_47 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_48 ),
    .SUM(tdc_inst_dl_capt_D_47 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_48_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_48 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_48 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_48 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_49 ),
    .SUM(tdc_inst_dl_capt_D_48 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_49_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_49 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_49 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_49 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_50 ),
    .SUM(tdc_inst_dl_capt_D_49 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_4_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_4 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_4 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_4 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_5 ),
    .SUM(tdc_inst_dl_capt_D_4 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_50_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_50 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_50 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_50 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_51 ),
    .SUM(tdc_inst_dl_capt_D_50 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_51_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_51 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_51 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_51 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_52 ),
    .SUM(tdc_inst_dl_capt_D_51 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_52_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_52 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_52 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_52 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_53 ),
    .SUM(tdc_inst_dl_capt_D_52 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_53_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_53 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_53 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_53 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_54 ),
    .SUM(tdc_inst_dl_capt_D_53 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_54_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_54 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_54 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_54 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_55 ),
    .SUM(tdc_inst_dl_capt_D_54 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_55_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_55 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_55 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_55 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_56 ),
    .SUM(tdc_inst_dl_capt_D_55 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_56_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_56 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_56 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_56 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_57 ),
    .SUM(tdc_inst_dl_capt_D_56 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_57_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_57 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_57 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_57 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_58 ),
    .SUM(tdc_inst_dl_capt_D_57 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_58_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_58 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_58 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_58 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_59 ),
    .SUM(tdc_inst_dl_capt_D_58 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_59_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_59 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_59 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_59 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_60 ),
    .SUM(tdc_inst_dl_capt_D_59 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_5_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_5 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_5 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_5 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_6 ),
    .SUM(tdc_inst_dl_capt_D_5 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_60_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_60 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_60 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_60 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_61 ),
    .SUM(tdc_inst_dl_capt_D_60 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_61_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_61 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_61 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_61 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_62 ),
    .SUM(tdc_inst_dl_capt_D_61 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_62_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_62 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_62 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_62 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_63 ),
    .SUM(tdc_inst_dl_capt_D_62 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_63_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_63 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_63 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_63 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_64 ),
    .SUM(tdc_inst_dl_capt_D_63 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_6_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_6 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_6 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_6 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_7 ),
    .SUM(tdc_inst_dl_capt_D_6 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_7_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_7 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_7 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_7 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_8 ),
    .SUM(tdc_inst_dl_capt_D_7 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_8_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_8 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_8 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_8 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_9 ),
    .SUM(tdc_inst_dl_capt_D_8 ));
 sky130_fd_sc_hd__fa_2 tdc_inst_dl_inst_dl_genblk_dl_rca_genblk_9_FA  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_9 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_b_int_9 ),
    .CIN(tdc_inst_dl_inst_dl_genblk_dl_c_9 ),
    .COUT(tdc_inst_dl_inst_dl_genblk_dl_c_10 ),
    .SUM(tdc_inst_dl_capt_D_9 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_0_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_0 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_10_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_10 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_11_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_11 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_12_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_12 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_13_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_13 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_14_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_14 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_15_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_15 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_16_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_16 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_17_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_17 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_18_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_18 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_19_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_19 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_1_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_1 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_20_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_20 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_21_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_21 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_22_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_22 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_23_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_23 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_24_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_24 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_25_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_25 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_26_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_26 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_27_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_27 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_28_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_28 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_29_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_29 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_2_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_2 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_30_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_30 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_31_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_31 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_32_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_32 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_33_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_33 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_34_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_34 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_35_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_35 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_36_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_36 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_37_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_37 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_38_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_38 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_39_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_39 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_3_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_3 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_40_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_40 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_41_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_41 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_42_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_42 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_43_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_43 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_44_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_44 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_45_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_45 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_46_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_46 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_47_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_47 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_48_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_48 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_49_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_49 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_4_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_4 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_50_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_50 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_51_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_51 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_52_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_52 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_53_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_53 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_54_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_54 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_55_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_55 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_56_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_56 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_57_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_57 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_58_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_58 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_59_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_59 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_5_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_5 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_60_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_60 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_61_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_61 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_62_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_62 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_63_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_63 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_6_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_6 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_7_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_7 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_8_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_8 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_zeros_const_zeros_genblk_9_const_zero  (.LO(tdc_inst_dl_inst_dl_genblk_dl_b_int_9 ));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_25 (.HI(net25));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_26 (.HI(net26));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_27 (.HI(net27));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_28 (.HI(net28));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_29 (.HI(net29));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_30 (.HI(net30));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_31 (.HI(net31));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_32 (.HI(net32));
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

