VERSION 1.0;

END LIBRARY
